-- Created on: 2000-09-04
-- Created by: Vincent DELOS
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Explorer from XBooleanOperations 

	---Purpose:  the explorer associated  to the Data Structure to
	--          retrieve   subshapes of a  given   shape stored in
	--          ShapesDataStructure.

uses
    Shape    from TopoDS,
    ShapeEnum from TopAbs,
    ShapesDataStructure from XBooleanOperations,
    PShapesDataStructure from XBooleanOperations

is
    Create (SDS: ShapesDataStructure)  
    	returns Explorer from XBooleanOperations;

    --modified by NIZNHY-PKV Sun Dec 15 16:24:39 2002  f 
    Delete(me:  out)  
    	is virtual; 
    ---C++:  alias  "Standard_EXPORT virtual ~XBooleanOperations_Explorer()  {Delete();}" 
    --modified by NIZNHY-PKV Sun Dec 15 16:27:53 2002  t 
    
    Init (me:in out;  
    	aShape: Integer;  
    	TargetToFind: ShapeEnum;  
    	TargetToAvoid: ShapeEnum = TopAbs_SHAPE) is virtual;
    
    Next (me:in out)  
    	is virtual;
    
    More (me)  
    	returns Boolean;
    
    Current (me:in out)  
    	returns Integer is virtual;

    Dump (me; S : in out OStream)  
    	is virtual;


fields

myShapesDataStructure: PShapesDataStructure is protected;
---Purpose: the data structure we're working on.

myStack : Address is protected;
---Purpose: contains all the numbers associated to the shapes.
myTopOfStack : Integer is protected;
---Purpose: gives the position of  the  highest element in the stack,
--          i.e. the index of the number of the current shape.
mySizeOfStack : Integer is protected;
---Purpose: gives the number of elements in the stack.

myTargetToFind : ShapeEnum is protected;
---Purpose: the kind of shape we are looking for.
myTargetToAvoid: ShapeEnum is protected;
---Purpose: the kind of shape we want to avoid.

hasMore : Boolean is protected;
---Purpose: if we still have a new shape to return.

end Explorer;
