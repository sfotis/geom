-- Created on: 2000-11-23
-- Created by: Michael KLOKOV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class Curve from XIntTools


uses
    Curve from Geom,
    Curve from Geom2d,
    Pnt  from gp, 
    CurveType from GeomAbs
is
    Create  
    	returns Curve from XIntTools;
	---Purpose:
	--- Empty constructor
	---

    Create(Curve3d: Curve from Geom;  
    	   FirstCurve2d : Curve from Geom2d;
    	   SecondCurve2d: Curve from Geom2d)
    	returns Curve from XIntTools;
	---Purpose:
	--- Initializes me by a 3d curve
	--- and two 2d curves
	---

    SetCurves(me: in out;  
    	      Curve3d: Curve from Geom;  
    	      FirstCurve2d  : Curve from Geom2d;
    	      SecondCurve2d : Curve from Geom2d);
    	---Purpose:
	--- Modifier
	---
    
    SetCurve(me: in out;  
    	    	Curve3d: Curve from Geom);
    	---C++: inline
	---Purpose:
	--- Modifier
	---
    
    SetFirstCurve2d(me: in out;  
    	    	FirstCurve2d: Curve from Geom2d);
    	---C++: inline
	---Purpose:
	--- Modifier
	---
    
    SetSecondCurve2d(me: in out;  
    	    	SecondCurve2d: Curve from Geom2d);
    	---C++: inline
	---Purpose:
	--- Modifier
	---

    Curve(me)  
    	returns any Curve from Geom;
    	---C++: return const &
	---C++: inline
	---Purpose:
	--- Selector
	---
    
    FirstCurve2d(me)
    	returns any Curve from Geom2d;
    	---C++: return const &
	---C++: inline
	---Purpose:
	--- Selector
	---
	    
    SecondCurve2d(me)
    	returns any Curve from Geom2d;
    	---C++: return const &
	---C++: inline 
	---Purpose:
	--- Selector
	---
	
    HasBounds (me) 
    	returns Boolean from Standard;
	---Purpose:
	--- Returns true if 3d curve is BoundedCurve from Geom
	---

    Bounds    (me; aT1:out Real from Standard;    	  
                   aT2:out Real from Standard;    	  
		   aP1:out Pnt  from gp;     
		   aP2:out Pnt  from gp);
    	---Purpose:
	--- Returns boundary parameters
	--- and corresponded 3d point.
	---
	--  Warning:
	--- If HasBounds returns false
	--- the returned parameters are equal
	--- to zero.
	---

    D0        (me;  
    	       aT1:out Real from Standard; 
               aP1:out Pnt  from gp) 
    	returns Boolean from Standard;
	---Purpose:
	--- Computes 3d point corresponded to parameter aT1
	--- Returns true if given parameter aT1
	--- is inside the boundaries of the curve
	---
     
    Type  (me) 
    	returns CurveType from GeomAbs; 
	---Purpose:
	--- Returns the type of 3d curve
	---
 
fields

    my3dCurve : Curve from Geom;
    my2dCurve1: Curve from Geom2d;
    my2dCurve2: Curve from Geom2d;
    
end Curve from XIntTools;
