-- Created on: 2001-02-08
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PaveFiller from XBOPTools 

	---Purpose:  The algorithm that provides  
        ---  1. creation of the data structure (DS)    	 
        ---  2. creation of the interferences' pool   	 
        ---  3. invocation of Perform() to fill the DS 
    	---   
        ---
uses
    
    PShapesDataStructure    from XBooleanOperations, 
    
    InterferencePool        from XBOPTools,  
    PInterferencePool       from XBOPTools,  
    PavePool                from XBOPTools, 
    CommonBlockPool         from XBOPTools, 
    SplitShapesPool         from XBOPTools, 
    
    Pave                    from XBOPTools,  
    PaveBlock               from XBOPTools,  
    PaveSet                 from XBOPTools, 
    Curve                   from XBOPTools,
    SSInterference          from XBOPTools, 
    ListOfPaveBlock         from XBOPTools, 
    IteratorOfCoupleOfShape from XBOPTools, 
    SSInterference          from XBOPTools, 
    SSIntersectionAttribute from XBOPTools, 
    ShrunkRange             from XIntTools, 
    Context                 from XIntTools, 
    
    ShapeEnum           from  TopAbs, 
    ListOfInteger       from TColStd, 
    IndexedMapOfInteger from TColStd, 
    
    Pnt     from gp,
    Vertex  from TopoDS,
    SetOfInteger  from  TColStd


is 
 
    Create   
    	returns PaveFiller from XBOPTools; 
    	---Purpose:  
    	--- Empty Contructor  
    	---
    Create  (aIP: InterferencePool from XBOPTools) 
    	returns PaveFiller from XBOPTools; 
    	---Purpose:   
    	--- Constructor 
    	---
    Create  (theIP              : InterferencePool from XBOPTools;
    	     theSectionAttribute: SSIntersectionAttribute from XBOPTools) 
    	returns PaveFiller from XBOPTools; 
    	---Purpose:   
    	--- Constructor
    	---
    Destroy (me: in out) 
	is  virtual;     
    	---C++: alias "Standard_EXPORT virtual ~XBOPTools_PaveFiller(){Destroy();}"     
    	---Purpose:   
    	--- Destructor
    	---
    Perform    (me:out) 
	is virtual;       
    	---Purpose:
    	--- Fills the DS               
    	---
 
    PartialPerform(me:out; anObjSubSet, aToolSubSet:  SetOfInteger  from  TColStd) 
	is virtual;       
       
    ToCompletePerform(me:out)		   
	is virtual;       
 
    PerformVV  (me:out) 
    	is  virtual protected; 
    	---Purpose:
    	--- Computes Vertex/Vertex interferences                
    	---
    PerformVE  (me:out) 
    	is  virtual protected;  
    	---Purpose:
    	--- Computes Vertex/Edge interferences                
    	---
    PerformVF  (me:out) 
    	is  virtual protected;  
    	---Purpose:
    	--- Computes Vertex/Face interferences                
    	---
    PerformEE  (me:out) 
    	is  virtual protected;  
    	---Purpose:
    	--- Computes Edge/Edge interferences                
    	---
    PerformEF  (me:out) 
    	is  virtual protected; 
    	---Purpose:
    	--- Computes Edge/Face interferences                
    	---
    PerformFF  (me:out) 
    	is  virtual protected;   
    	---Purpose:
    	--- Computes Face/Face interferences                
    	---

    -------------------------------------------------------------- 
    --- 
    ---	  Selectors   
    ---   
    --- 
    SetContext(me:out; 
    	    aContext:  Context from XIntTools); 
    	---Purpose:
    	--- Sets the intersecton context                 
    	---   
    Context(me) 
    	 returns Context from XIntTools; 
    	---C++:return const &	
    	---Purpose:
    	--- Selector                
    	---
--    ChangeContext(me:out) 
--    	 returns Context from XIntTools;  
    	--  C++:return &	
    	---Purpose:
    	--- Selector                
    	---
    SetInterferencePool(me:out; 
    	 aPool:InterferencePool from XBOPTools); 
    	---Purpose:
    	--- Selector                
    	---
    IsDone(me) 
    	returns  Boolean  from  Standard;  
    	---Purpose:
    	--- Selector
    	---
    PavePool(me) 
    	returns  PavePool from XBOPTools; 
    	---C++:return const &	 
    	---Purpose:
    	--- Selector               
    	---
    ChangePavePool(me:out) 
    	returns  PavePool from XBOPTools; 
    	---C++:return &	
   	---Purpose:
    	--- Selector               
    	---
    CommonBlockPool(me) 
    	returns  CommonBlockPool from XBOPTools; 
    	---C++:return const &	 
    	---Purpose:
    	--- Selector               
    	---
    ChangeCommonBlockPool(me:out) 
    	returns  CommonBlockPool from XBOPTools; 
    	---C++:return &	
    	---Purpose:
    	--- Selector               
    	---
    SplitShapesPool(me)  
    	returns  SplitShapesPool from XBOPTools;
    	---C++:return const &	
    	---Purpose:
    	--- Selector               
    	---

    ChangeSplitShapesPool(me:out)  
    	returns  SplitShapesPool from XBOPTools;
    	---C++:return  &	
    	---Purpose:
    	--- Selector               
    	---
    DS(me:out) 
    	returns PShapesDataStructure from XBooleanOperations;  
    	---Purpose:
    	--- Selector               
    	---
    InterfPool(me:out) 
    	returns PInterferencePool from XBOPTools; 
    	---Purpose:
    	--- Selector               
    	---
 
    IteratorOfCoupleOfShape(me)  
    	returns  IteratorOfCoupleOfShape from XBOPTools;
    	---C++:return const &	
    	---Purpose:
    	--- Selector               
	---
      
    SectionAttribute(me)
    	returns SSIntersectionAttribute from XBOPTools;
    	---C++: return const &
    	---Purpose:
    	--- Selector   
	---

    SetSectionAttribute(me:out; 
    	anAtt  :  SSIntersectionAttribute from XBOPTools);
    	---Purpose:
    	--- Selector       
	---
    -------------------------------------------------------------- 
    ---	     
    ---  PaveBlocks for Split Parts of Edges.  
    ---     
    --- 
    SortTypes      (me;   
    	    anInd1:in out Integer from Standard; 
            anInd2:in out Integer from Standard) 
    	is protected;  
    	---Purpose:
    	--- Sorts the types of shapes with DS-indices  
    	--- <anInd1> and  <anInd2> in increasing order of  
    	--- types of the shapes               
    	---
    PerformNewVertices  (me:out) 
    	is protected;     	     
     
    IsSuccesstorsComputed (me;  
    	    iF1:Integer from  Standard; 
    	    iF2:Integer from  Standard) 
    	returns  Boolean from Standard 
    	is protected;    
     
    PrepareEdges  (me:out) 
    	is virtual protected;  
    	---Purpose:   
    	--- Prepare end paves for each edge 
    	---
    PreparePaveBlocks (me:out; 
    	    	    	aType1: ShapeEnum  from  TopAbs; 
    	    	    	aType2: ShapeEnum  from  TopAbs) 
    	is virtual protected; 
    	---Purpose:   
    	--- Prepare PaveBlocks  for  each  edge  (EE-interferences) 
    	---
    PreparePaveBlocks (me:out;   
    	    	       anE:Integer from Standard) 
    	is virtual protected;  
    	---Purpose:  
    	--- Prepare PaveBlocks for given edge (EE-interferences) 
    	---
    RefinePavePool(me:out) 
    	is protected;  
    	---Purpose:  
    	--- Refines myPavePool taking into account new Paves obtained from EE algo 
    	---
    MakeSplitEdges(me:out) 
    	is protected;   
    	---Purpose:  
    	--- Makes split edges from source edges 
    	---
    DoSDEdges(me:out) 
    	is protected;    
    	---Purpose:
    	--- Update Lists of PaveBlocks with info about 
    	--- indices of split edges that are Same Domain 
    	--- with other splits or faces 
    	---
    CorrectShrunkRanges(me:out; 
    	    	    	aSide:  Integer  from  Standard; 
    	    	    	aPave:  Pave from XBOPTools; 
    	    	    	aSR  :  out ShrunkRange  from  XIntTools)
    	is protected;  
    	---Purpose:
    	--- Update Shrunk  Range <aSR> for Pave <aPave> 
    	---
    SplitIndex  (me:out;  aPB:PaveBlock from XBOPTools)  
    	returns Integer from Standard 
    	is protected;  
    	---Purpose:  
    	--- Returns  the Index of Split edge for the PaveBlock <aPB> 
    	--- in  DS. 
    	--- If the PaveBlock is not found, returns 0; 
    	---
    IsBlocksCoinside (me; 
    	aPB1:PaveBlock from XBOPTools;
    	aPB2:PaveBlock from XBOPTools) 
	returns Boolean from Standard 
    	is protected;   
    	---Purpose: 	 
    	--- Returns  TRUE if the two PaveBlocks have vertices 
    	--- that touch each other in terms of Tolerances of 
    	--- the vertices 	     
    	---
    -------------------------------------------------------------- 
    ---	  
    ---  Some of API FUNCTIONS  
    --- 
    --- 
    SplitsInFace(me:out; 
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the face <nF1> get all splits that are IN-2D          
    	--- to  the face <nF2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
    SplitsInFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the edge <nE1> get all splits that are IN-2D          
    	--- to  the face <nF1>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
    SplitsOnEdge(me:out; 
    	         nE1 :Integer from Standard;  
    	         nE2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the edge <nE1> get all splits that are ON-3D          
    	--- to  the edge <nE2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
    SplitsOnFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the edge <nE1> get all splits that are ON-3D          
    	--- to  the face <nF2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
    SplitsOnFace(me:out;  
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfInteger from TColStd) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the face <nF1> get all splits that are ON-3D          
    	--- to  the face <nF2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
     
    SplitsInFace(me:out; 
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from XBOPTools) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the face <nF1> get all PaveBlocks that are IN-2D          
    	--- to  the face <nF2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
     
    SplitsInFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from XBOPTools) 
    	returns Integer from Standard;  
    	---Purpose:   
    	--- For the edge <nE1> get all PaveBlocks that are IN-2D          
    	--- to  the face <nF1>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
     
    SplitsOnEdge(me:out; 
    	         nE1 :Integer from Standard;  
    	         nE2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from XBOPTools) 
    	returns Integer from Standard;  
    	---Purpose:   
    	--- For the edge <nE1> get all PaveBlocks that are ON-3D          
    	--- to  the edge <nE2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
     
    SplitsOnFace(me:out; 
    	         nE1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from XBOPTools) 
    	returns Integer from Standard;  
    	---Purpose:  
    	--- For the edge <nE1> get all PaveBlocks that are ON-3D          
    	--- to  the face <nF2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---

    SplitsOnFace(me:out;  
    	         aBid:Integer from Standard;  
    	         nF1 :Integer from Standard;  
    	         nF2 :Integer from Standard;  
    	         aLs :out ListOfPaveBlock from XBOPTools) 
    	returns Integer from Standard;  
    	---Purpose: 
    	--- For the face <nF1> get all PaveBlocks that are ON-3D          
    	--- to  the face <nF2>; The result is in <aLs> 
    	--- Returns 0 if OK; 
    	---
    FindSDVertex (me; 
    	    	    nV:  Integer  from  Standard) 
    	returns Integer from Standard; 
    	---Purpose:
    	--- Find  for the vertex <nV> SD-vertex (if possible) and return  
    	--- its DS-index.  Otherwise it returns 0.
	---
     
    --------------------------------------------------------------- 
    ---	  
    ---   Section  Edges.  Protected Block.
    --- 
    ---	     
    MakeBlocks(me:out) 
    	is protected; 
    	---Purpose: 
    	--- Make Pave Blocks for intersection curves    
    	---
    MakeAloneVertices(me:out) 
    	is protected; 
    	---Purpose: 
    	--- Make vertices that are place of intersection  
    	--- between faces       
    	---
    PutPaveOnCurve(me:out; 
    	    	   aPaveSet: PaveSet from XBOPTools; 
		   aTolR3D : Real from Standard; 				   		     
    	    	   aBCurve :out Curve from XBOPTools) 
       	is protected;   
    	---Purpose: 
    	--- Among Paves from <aPaveSet> find ones that belong 
    	--- to intersection curve <aBCurve> with 3D-tolerance  
    	--- value <aTolR3D>
    	---
    PutPaveOnCurve(me:out; 
    	    	   aPave   : Pave from XBOPTools; 
    	    	   aTolR3D : Real from Standard;  
    	    	   aBCurve :out Curve from XBOPTools) 
       	is protected;     
    	---Purpose: 
    	--- Try to put Pave <aPave> on intersection curve <aBCurve>  
    	--- with 3D-tolerance value <aTolR3D>
    	---

    PutPavesOnCurves(me:out)
    	is protected;

    PrepareSetForFace(me:out;  
    	    	    nF1 :Integer from Standard;  
    	    	    nF2 :Integer from Standard;  
	    	    aPaveSet:out PaveSet from XBOPTools); 
    	---Purpose:  
    	--- For couple of faces <nF1>, <nF2> prepare set of all paves 
    	--- of all edges <aPaveSet>
    	---
    MakeSectionEdges(me:out) 
    	is protected;  
    	---Purpose:  
    	--- For all inrefered faces make section edges from  
    	--- intersection curves and corresp.  Paves on them      
    	---
    PutBoundPaveOnCurve (me:out; 
    	    	    aBC :out Curve from XBOPTools;	 
     	    	    aFF :out SSInterference from XBOPTools) 
    	is protected; 
    	---Purpose: 	     
    	--- Try to  put own  bounds of the curve on the curve <aBC> 
    	---
    PutBoundPaveOnCurve (me:out;  
    	    	    aP  : Pnt from  gp; 
		    aT  : Real from Standard; 			 
    	    	    aBC :out Curve from XBOPTools;	 
     	    	    aFF :out SSInterference from XBOPTools) 
    	is protected;  
    	---Purpose: 	     
    	--- Try to put 3D-point <aP> (parameter aT)  on the curve <aBC> 
    	---
    PutBoundPaveOnCurveSpec (me:out; 
    	    	    aBC :out Curve from XBOPTools;	 
     	    	    aFF :out SSInterference from XBOPTools) 
    	is protected; 
    	---Purpose: 	     
    	--- Try to  put own  bounds of the curve on the curve <aBC> 
    	--- 
    PutBoundPaveOnCurveSpec (me:out;  
    	    	    aP  : Pnt from  gp; 
		    aT  : Real from Standard; 			 
    	    	    aBC :out Curve from XBOPTools;	 
     	    	    aFF :out SSInterference from XBOPTools) 
    	is protected;  
    	---Purpose: 	     
    	--- Try to put 3D-point <aP> (parameter aT)  on the curve <aBC> 
    	--- 
 
--modified by NIZNHY-PKV Thu Oct 20 07:17:11 2011f 
    PutClosingPaveOnCurve (me:out; 
    	    	    aBC :out Curve from XBOPTools;	 
     	    	    aFF :out SSInterference from XBOPTools)  
	is protected; 
	---Purpose: 	     
    	--- Put paves on the curve <aBC> in case when <aBC>   
        --  is closed 3D-curve  
    	---      
--modified by NIZNHY-PKV Thu Oct 20 07:17:11 2011t	 

    FindPave            (me:out; 
		    aP  :Pnt from  gp;  
    	    	    aTpV: Real from Standard;  
    	    	    aPS: PaveSet from XBOPTools; 
		    aPV:out Pave from XBOPTools) 
    	returns Boolean from Standard
       	is protected; 
    	---Purpose: 	     
    	--- Returns TRUE if 3D-point <aP> coinsides with some Pave 
    	--- from <aPS> (with 3D-tolerance value <aTpV>); 
    	--- In  TRUE case <aPV> will contain the Pave  .      	     
    	---
    CheckCoincidence(me:out;  
    	    	    aPB: PaveBlock      from XBOPTools;  
     	    	    aFF: SSInterference from XBOPTools) 
    	returns Boolean from Standard 
    	is protected;  
    	---Purpose: 	     
    	--- Returns TRUE if PaveBlock <aPB> lays on the faces 
    	--- from FF-interference <aFF> 
    	---
    CheckIntermediatePoint(me:out;  
    	    	    aPB : PaveBlock      from XBOPTools;  
    	    	    aPBR: PaveBlock      from XBOPTools;  
     	    	    aTol: Real  from  Standard) 
    	returns Integer from Standard 
    	is protected;  
    	---Purpose: 	     
    	--- Returns 0 if some arbitrary intermediate point from   
    	--- PaveBlock <aPB> lays on the PaveBlock  <aPBR> 
    	--- (with 3D-tolerance value <aTol>)
    	---
 
    CheckFacePaves(me:out;  
    	    	    aV : Vertex  from TopoDS;  
     	    	    nF:  Integer from Standard) 
    	returns Integer from Standard 
    	is protected; 
    	---Purpose: 	 
    	--- Internal  usage 
    	---
    StickVertices (me:out;   
    	    	    nF1:  Integer from Standard;
    	    	    nF2:  Integer from Standard; 
		    aMV:out IndexedMapOfInteger from TColStd) 
	is protected; 	    
    	---Purpose: 	 
    	--- Internal  usage 
    	---
    ExpectedPoolLength(me) 
    	returns  Integer from Standard 
	is protected;
    	---Purpose: 	 
    	--- Returns the value of expected length of array of interferences 
    	---

    RestrictCurveIn2d(me: in out; nE, nF1, nF2    : Integer from Standard;
    	    			theTolerance: Real from Standard;
			     	theBC       : in out Curve from XBOPTools)
    	is private;

    RecomputeCommonBlocks(me: in out; nE: Integer from Standard)
    	is private;

    ExtendedTolerance(me:out; 
    	    nV      : Integer from Standard; 
            aTolExt : out Real from Standard) 
	returns Boolean from Standard 		     
	is  protected;		     

fields 
 
    myIntrPool         :  PInterferencePool from XBOPTools
    	is protected;
    myDS               :  PShapesDataStructure from XBooleanOperations 
    	is protected;   
    myPavePool         :  PavePool from XBOPTools 
    	is protected; 
    myPavePoolNew      :  PavePool from XBOPTools 
    	is protected; 
    myCommonBlockPool  :  CommonBlockPool from XBOPTools 
    	is protected;  
    mySplitShapesPool  :  SplitShapesPool from XBOPTools 
    	is protected; 
    mySectionAttribute :  SSIntersectionAttribute from XBOPTools 
    	is protected;
    myNbSources        :  Integer from Standard 
    	is protected; 
    myNbEdges          :  Integer from Standard 
    	is protected;      
    myIsDone           :  Boolean from Standard 
    	is protected; 
    myDSIt             :  IteratorOfCoupleOfShape from XBOPTools 
    	is protected; 
    myContext           :  Context from XIntTools 
    	is protected;  	     

end PaveFiller;
