-- Created on: 2000-11-22
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


package XBOPTColStd 
     
    ---Purpose: 
     ---         Contains auxiliary classes used  by   
    ---          boolean  operations algorithm.  
    
uses  
    gp,   
    TopoDS,  
    TopTools,
    TCollection, 
    TColStd  
---
is    

    generic class CArray1;
    ---Purpose:  
    --  The class represents unidimensionnal arrays
    --  of fixed size known at run time.  
    --  Run-time boundary check is performed
    --  The range of the index is user defined from 0 to Length-1 
    --
    class  Dump; 
    --  The class provides dump service used for debugging   
    --  purposes 
    --  
    class Failure;       
    --  The class provides exception objects 
    --  
    class ShapeWithRank;         	 
    --  The auxiliary class provides structure to store a shape 
    --  and its rank 
    ---     
    class ShapeWithRankHasher; 
    --  The auxiliary class provides hash code for mapping 
    --  ShapeWithRank objects 
    ---   
    ---
    ---                 I  n  s  t  a  n  t  i  a  t  i  o  n  s  
    ---       
    class  CArray1OfInteger  instantiates  
    	CArray1 from XBOPTColStd(Integer from Standard);  
	 
    class CArray1OfShape instantiates  
    	CArray1 from XBOPTColStd(Shape from TopoDS);  
	 
    class CArray1OfPnt2d instantiates  
    	CArray1 from XBOPTColStd(Pnt2d from gp);   
     
    class  IndexedDataMapOfIntegerInteger  instantiates 
    	IndexedDataMap from TCollection  (Integer, 
	    	    	    	    	  Integer,  
	    	    	    	    	  MapIntegerHasher from TColStd);  
    class  ListOfListOfShape instantiates 
    	List from TCollection (ListOfShape from TopTools);

    class  IndexedDataMapOfIntegerIndexedMapOfInteger  instantiates 
    	IndexedDataMap from TCollection  (Integer, 
	    	    	    	    	  IndexedMapOfInteger from TColStd,    
	    	    	    	    	  MapIntegerHasher from TColStd); 

    class  IndexedDataMapOfSWRInteger instantiates 
    	IndexedDataMap from TCollection  (ShapeWithRank, 
	    	    	    	    	  Integer from Standard,    
	    	    	    	    	  ShapeWithRankHasher from XBOPTColStd);
    
    
     

end  XBOPTColStd;
