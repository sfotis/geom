-- Created on: 2001-08-02
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class FaceInfo from XBOP 

	---Purpose: 
    	---  The  auxiliary class to store data about faces on a  shell 
    	---  that have common edge         	 
	---  
	
uses
    Face  from TopoDS, 
    Pnt   from gp, 
    Dir   from gp,
    Pnt2d from gp 
    
--raises

is 
    Create 
    	returns FaceInfo from XBOP;
    	---Purpose:  
    	--- Empty constructor;  
    	---
    SetFace   (me:out; 
    	        aF:Face from TopoDS); 
    	---Purpose: 
    	--- Modifier
    	---
    SetPassed (me:out;   
    	        aFlag:Boolean from Standard); 
    	---Purpose: 
    	--- Modifier
    	---
    SetPOnEdge (me:out;   
    	        aP:Pnt from gp);  
    	---Purpose: 
    	--- Modifier
    	---
    SetPInFace (me:out;   
    	        aP:Pnt from gp);   
    	---Purpose: 
    	--- Modifier
    	---
    SetPInFace2D (me:out;   
    	        aP:Pnt2d from gp);
    	---Purpose: 
    	--- Modifier
    	---
    SetNormal (me:out;   
    	        aD:Dir from gp);   
    	---Purpose: 
    	--- Modifier
    	---
    SetAngle  (me:out;   
    	        A:Real from Standard); 
    	---Purpose: 
    	--- Modifier
    	---
     
    Face      (me) 
    	returns Face from TopoDS; 
    	---C++:  return const & 
    	---Purpose: 
    	--- Selector
    	---
    POnEdge   (me) 
	returns Pnt from gp; 
    	---C++:  return const &  
    	---Purpose: 
    	--- Selector
    	---
    PInFace   (me) 
	returns Pnt from gp; 
    	---C++:  return const &  
    	---Purpose: 
    	--- Selector
    	---
    PInFace2D   (me) 
	returns Pnt2d from gp; 
    	---C++:  return const &  
    	---Purpose: 
    	--- Selector
    	---
 
    Normal   (me) 
	returns Dir from gp; 
    	---C++:  return const &  
    	---Purpose: 
    	--- Selector
    	---
    IsPassed (me)   
    	returns Boolean from Standard; 
    	---Purpose: 
    	--- Selector
    	---
    Angle  (me)   
    	returns Real from Standard; 
    	---Purpose: 
    	--- Selector
    	---
fields  

    myFace  : Face from TopoDS; 
    myPassed: Boolean from Standard; 
    myPOnEdge  :  Pnt from gp;  
    myPInFace  :  Pnt from gp; 
    myPInFace2D:  Pnt2d from gp; 
    myNormal   :  Dir from gp;  
    myAngle    :  Real from  Standard; 

end FaceInfo;
