-- Created on: 2000-09-07
-- Created by: Vincent DELOS
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class OnceExplorer from XBooleanOperations  
    inherits Explorer from XBooleanOperations

	---Purpose: 

uses
    Shape     from TopoDS,
    ShapeEnum from TopAbs,
    ShapesDataStructure from XBooleanOperations,
    PShapesDataStructure from XBooleanOperations

--raises

is
    Create (SDS: ShapesDataStructure)  
    	returns OnceExplorer from XBooleanOperations;
--modified by NIZNHY-PKV Sun Dec 15 16:24:39 2002  f 
    Delete(me:  out)  
    	is redefined virtual; 
    ---C++:  alias  "Standard_EXPORT virtual ~XBooleanOperations_OnceExplorer()  {Delete();}"
--modified by NIZNHY-PKV Sun Dec 15 16:24:42 2002  t
    
    Init (me:in out;  
    	    aShape: Integer;  
    	    TargetToFind: ShapeEnum;  
    	    TargetToAvoid: ShapeEnum = TopAbs_SHAPE) is redefined;
    
    Next (me:in out)  
    	is redefined;
    	
    Current (me:in out)  
    	returns Integer is redefined;

    Dump (me; S : in out OStream)  
    	is redefined; 


fields

    myArrayOfBits : Address;
    ---Purpose: to say if we already visited a shape.
    mySizeOfArrayOfBits : Integer;
    ---Purpose: the size of <myArrayOfBits>.

end OnceExplorer;
