-- Created on: 2001-12-13
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PntOn2Faces from XIntTools 

	---Purpose: Contains two points PntOnFace from XIntTools and a flag

uses
    PntOnFace from XIntTools
---raises

is 
    Create 
    	returns PntOn2Faces from XIntTools; 
	---Purpose:
	--- Empty constructor
	---
	 
    Create(aP1:	PntOnFace from XIntTools;
           aP2:	PntOnFace from XIntTools);
    	---Purpose:
	--- Initializes me by two points aP1 and aP2
	---
	    
    SetP1 (me:out; 
    	aP1: PntOnFace from XIntTools);
	---Purpose:
	--- Modifier
	---
	 
    SetP2 (me:out; 
    	aP2: PntOnFace from XIntTools);
	---Purpose:
	--- Modifier
	---

    SetValid(me:out; 
	bF : Boolean from Standard); 
	---Purpose:
	--- Modifier
	---
     
    P1(me) 
    	returns PntOnFace from XIntTools; 
    	---C++:  return const &  
	---Purpose:
	--- Selector
	---
     
    P2(me) 
    	returns PntOnFace from XIntTools; 
    	---C++:  return const & 
	---Purpose:
	--- Selector
	---

    IsValid(me) 
	returns Boolean from Standard; 
	---Purpose:
	--- Selector
	---

fields
  
    myIsValid : Boolean from Standard;    
    myPnt1    : PntOnFace from XIntTools;
    myPnt2    : PntOnFace from XIntTools;
    
     
end PntOn2Faces;
