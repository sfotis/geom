-- Created on: 2001-05-31
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Draw from XBOP 

	---Purpose: 
    	---  auxiliary class to display intermediate results  
    	---  in  Draw's winowds for the debugging purposes 
	---   
	 
uses
    ListOfShape from TopTools,
    Face from TopoDS,
    Edge from TopoDS 
    
is
    DrawListOfShape  (myclass; 
    	aList  : ListOfShape from TopTools; 
	aName  : CString from Standard); 
    	---Purpose:  
    	--- Display in  3D-view shapes from the ListOfShape  <aList>   
    	--- aName is base name of shape. Actual name for  each 
    	--- subsequent shape  will  be  aName+"_#",  where 
    	--- # - is ordered index of the shape in <aList>     	     
    	---
    DrawListOfEdgesWithPC  (myclass; 
	aFace  : Face from TopoDS;   		    		     
    	aList  : ListOfShape from TopTools; 
	aName  : CString from Standard);  
    	---Purpose:  
    	--- Display in  2D-view the edges from the ListOfShape  <aList>,  
    	--- that have P-curves for  the face <aFace>          
    	--- aName is base name of shape. Actual name for  each 
    	--- subsequent shape  will  be  aName+"_#",  where 
    	--- # -  is ordered index of the shape in <aList>     	     
    	---
    DrawListOfEdgesWithPC  (myclass; 
	aFace  : Face from TopoDS;   		    		     
    	aList  : ListOfShape from TopTools; 
	anInd  : Integer from Standard;         
    	aName  : CString from Standard);  
    	---Purpose:  
    	--- Display in  2D-view the edges from the ListOfShape  <aList>,  
    	--- that have P-curves for  the face <aFace>          
    	--- aName is base name of shape. Actual name for  each 
    	--- shape  will  be  aName+"_anInd"
	---
    DrawEdgeWithPC  (myclass; 
	aFace  : Face from TopoDS;   		    		     
    	aEdge  : Edge from TopoDS; 
	aName  : CString from Standard);   
    	---Purpose:   	
    	--- Display in  2D-view the edge,  
    	--- that has  P-curve for  the face <aFace>          
    	--- aName is the name of shape.  
    	---
    Wait(myclass); 
    	---Purpose:    
    	--- Wait  for  user's keystroke       
    	---
		    	    	
end Draw;
