-- Created on: 2000-11-27
-- Created by: Michael KLOKOV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class IteratorOfCoupleOfShape from XBOPTools

    	---Purpose: The class IteratorOfCoupleOfShape provides the iteration
    	---         on the couples of shapes stored in ShapesDataStructure 
	---         according to the given types of shapes and
	---         status of their intersection.
	---         The statuses are stored in 2 dimension array.

uses
    ShapeEnum from TopAbs,
    HArray2OfIntersectionStatus from XBOPTools,
    PShapesDataStructure from XBooleanOperations,
    IntersectionStatus from XBOPTools, 
    ListOfCoupleOfInteger from XBOPTools, 
    ListIteratorOfListOfCoupleOfInteger from XBOPTools,    
    NoSuchObject from Standard 
    
raises NoSuchObject from Standard 

is

    Create  
    	returns IteratorOfCoupleOfShape from XBOPTools;
    	---Purpose: 
    	--- Empty Constructor 
    	---

    Create(PDS: PShapesDataStructure from XBooleanOperations;
	   Type1: ShapeEnum from TopAbs;
    	   Type2: ShapeEnum from TopAbs)
    	returns IteratorOfCoupleOfShape from XBOPTools;
    	---Purpose: 
    	--- Initializes iterator by ShapesDataStructure and
    	--- shape types
	---

    Destroy(me: in out) is virtual;
        ---C++: alias "Standard_EXPORT virtual ~XBOPTools_IteratorOfCoupleOfShape(){Destroy();}"

    Initialize(me: in out; Type1: ShapeEnum from TopAbs;
    	    	    	   Type2: ShapeEnum from TopAbs) 
							    
	raises NoSuchObject from Standard 
    	is virtual;
    	---Purpose: 
    	--- Initializes iterator with shape types. 
    	--- The iterator uses PDS assigned in constructor or in SetDataStructure().
    	--- Raises the exception if myPDS is null.
	---


    SetDataStructure(me: in out; PDS: PShapesDataStructure from XBooleanOperations)
    	raises
	    NoSuchObject from Standard;
    	---Purpose: 
    	--- Initialize iterator with ShapeDataStructure.
	---
    

    More(me)  
    	returns Boolean from Standard 
    	is virtual;
	---Purpose:
	--- Returns True if there are still not
	--- treated couples of shapes
	---
    
    Next(me: in out) 
    	is virtual;
    	---Purpose:
	--- Moves to the next couple of iteration
	---
    
    Current(me; Index1: in out Integer from Standard;
    	    	Index2: in out Integer from Standard;
    	    	WithSubShape: out Boolean from Standard) 
    	is virtual;
    	---Purpose: 
    	--- Returns current couple of indices and
    	--- flag WithSubShape which is true 
    	--- if bounding boxes of subshapes
    	--- are intersected
	---

    ListOfCouple(me) 
    	returns  ListOfCoupleOfInteger from XBOPTools;  
    	---C++:  return const &
	---Purpose:
	--- Returns a list of couples of shape indices
	--- according to shape types by which
	--- the iterator was initialized
	---
	
    MoreP(me)  
    	returns Boolean from Standard   
    	is protected;
    
    NextP(me: in out) 
    	is protected;
    
    CurrentP(me;Index1: in out Integer from Standard;
    	    	Index2: in out Integer from Standard)
    	raises NoSuchObject from Standard 
    	is protected;

    SetIntersectionStatus(me: in out; Index1: Integer from Standard;
		        	      Index2: Integer from Standard;
    	    	    	    	      theStatus: IntersectionStatus from XBOPTools);
    	---Purpose:
	--- Sets status to array according to Index1 and Index2
	---

    GetTableOfIntersectionStatus(me)
    	returns HArray2OfIntersectionStatus from XBOPTools;
	---C++: return const &
	---Purpose:
	--- Returns 2 dimension array of intersection statuses
	---
    
    DumpTableOfIntersectionStatus(me);
    	---Purpose:
	--- For internal use
	---
    
fields
    myPDS: PShapesDataStructure from XBooleanOperations is protected;
    myTableOfStatus: HArray2OfIntersectionStatus from XBOPTools is protected;
    myCurrentIndex1: Integer from Standard is protected;
    myCurrentIndex2: Integer from Standard is protected;
    myType1:         ShapeEnum from TopAbs is protected;
    myType2:         ShapeEnum from TopAbs is protected;
--  
    myFirstLowerIndex :Integer from Standard is protected; 
    myFirstUpperIndex :Integer from Standard is protected; 
    mySecondLowerIndex:Integer from Standard is protected; 
    mySecondUpperIndex:Integer from Standard is protected; 
    myListOfCouple    :ListOfCoupleOfInteger from XBOPTools is protected;  
    myIterator        :ListIteratorOfListOfCoupleOfInteger from XBOPTools is protected;  
--  
end IteratorOfCoupleOfShape from XBOPTools;
