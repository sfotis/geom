-- Created on: 2000-05-18
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Range from XIntTools 

	---Purpose: The class describes the  1-d range 
        --          [myFirst, myLast].  	 

--uses
is 
    Create   
    	returns  Range from XIntTools ;
	---Purpose:
	--- Empty constructor
	---
     
    Create  (aFirst:Real  from  Standard;  aLast:Real  from  Standard) 
    	returns  Range from XIntTools ; 
	---Purpose:
	--- Initialize me by range boundaries
	---
	 
    SetFirst(me:out; aFirst:Real  from  Standard); 
    	---Purpose:
	--- Modifier
	---
     
    SetLast (me:out; aLast:Real  from  Standard);  
    	---Purpose:
	--- Modifier
	---
     
    First   (me) 
    	returns  Real  from  Standard; 
	---Purpose:
	--- Selector
	---
     
    Last   (me) 
    	returns  Real  from  Standard;  
	---Purpose:
	--- Selector
	---
	 
    Range  (me; aFirst:out Real  from  Standard;   
    	    	aLast :out Real  from  Standard);
    	---Purpose:
	--- Selector
	---
	    	
fields
    myFirst:  Real  from  Standard;
    myLast :  Real  from  Standard;
end Range;
