-- Created on: 2001-02-16
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ComparePave from XBOPTools 

	---Purpose: 
	---    	 
    	--- Auxiliary class for sorting paves along the edge    
        --- in acoordance with increasing order of parameter     
	    	 
uses 
    Pave from XBOPTools 
     
is
    Create   
    	returns ComparePave from XBOPTools; 
    	---Purpose:  
    	--- Empty constructor 
    	--- Default comparing tolerance value=1.e-12 
    	---
    Create  (aTol:Real from Standard) 
    	returns ComparePave from XBOPTools;  
    	---Purpose:   
    	--- Constructor that use comparing tolerance value as parameter.     
    	---
    IsLower (me; Left, Right: Pave from XBOPTools) 
    	returns Boolean ;
    	---Purpose:  
    	--- Returns True if <Left> is lower than <Right>. 
    	---
    IsGreater (me; Left, Right: Pave from XBOPTools) 
    	returns Boolean from Standard ;
    	---Purpose:  
    	--- Returns True if <Left> is greater than <Right>.
    	---
    IsEqual(me; Left, Right: Pave from XBOPTools) 
    	returns Boolean from Standard ; 
    	---Purpose:  
    	--- Returns True when <Right> and <Left> are equal.
    	---
	 
fields
    myTol: Real from Standard;  
     
end ComparePave;
