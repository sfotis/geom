-- Created on: 2002-02-04
-- Created by: Peter KURNEV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class StateFiller from XBOPTools 

	---Purpose:  
    	---  root class to compute states (3D)    
	---

uses 
    PaveFiller  from XBOPTools,
    PPaveFiller from XBOPTools, 
    PInterferencePool from XBOPTools, 
    PShapesDataStructure from XBooleanOperations, 
    
    Shape from TopoDS,   
    Edge  from TopoDS,
    State from TopAbs, 
    ShapeEnum from TopAbs,
    StateOfShape from XBooleanOperations
--raises

is 
    Create (aFiller: PaveFiller from XBOPTools) 
    	returns StateFiller from XBOPTools; 
    	---Purpose:  
    	--- Constructor 
    	---
    Do(me:out) 
    	is virtual; 
    	---Purpose: 
    	--- Launch the Filler   
    	---
    IsDone(me) 
    	returns Boolean from Standard; 
    	---Purpose:  
    	--- Returns true if Ok
	---
     
    ConvertState (myclass; 
    	    aSt: State from  TopAbs) 
	returns StateOfShape from XBooleanOperations; 
    	---Purpose:  
    	--- Convert conventional states to VDS-states
    	---
    ConvertState (myclass; 
    	    aSt: StateOfShape from XBooleanOperations) 
	returns State from  TopAbs; 
    	---Purpose:  
    	--- Convert VDS-states to conventional states     
    	---
    ClassifyEdgeToSolidByOnePoint  (me:out;  
    	    anEdge: Edge from TopoDS; 
	    aRef  : Shape from TopoDS)  
	returns State from  TopAbs;    
    	---Purpose:  
    	--- Computation the 3D-state of the edge <anEdge>  
    	--- to solid  <aRef>       
    	---
    ClassifyShapeByRef  (me:out; 
    	    aShape: Shape from TopoDS; 
    	    aRef  : Shape from TopoDS) 
    	returns  StateOfShape from XBooleanOperations;    
    	---Purpose:  
    	--- Computation the 3D-state of the shape <aShape>  
    	--- to solid <aRef>       
    	---
    SubType (myclass; 
    	    	aShape: Shape from TopoDS) 
    	returns ShapeEnum from TopAbs;    
    	---Purpose:  
    	--- Returns first subtype of <Shape> 
    	---
fields
    myFiller  : PPaveFiller from XBOPTools                    
    	is protected; 
    myDS      : PShapesDataStructure from XBooleanOperations  
    	is protected;   
    myIntrPool: PInterferencePool from XBOPTools              
    	is protected;  
    myIsDone  : Boolean   from Standard                      
    	is protected;  
     
end StateFiller;
