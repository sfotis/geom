-- Created on: 2001-02-08
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PaveSet from XBOPTools 

	---Purpose: 
    	-- class for storing/sorting paves that   
    	-- belong to an edge

uses
    ListOfPave from XBOPTools, 
    Pave       from XBOPTools

is 
    Create 
    	returns PaveSet from XBOPTools; 
    	---Purpose:  
    	--- Empty constructor 
    	---
    ChangeSet(me:out) 
    	returns ListOfPave from XBOPTools; 
    	---C++:  return & 
    	---Purpose:  
    	--- Access to the  list  
    	---
    Set(me) 
    	returns ListOfPave from XBOPTools; 
    	---C++:  return const & 	   
    	---Purpose:  
    	--- Access to the  list const 
    	---
    Append  (me:out; aPave:Pave from XBOPTools);
    	---Purpose:  
    	--- Appends <aPave>  to the  list  
    	---
    SortSet (me:out); 
    	---Purpose:  
    	--- Sorts  list in increasing order of paves' parameters 
    	---

fields 
    myPaveList: ListOfPave from XBOPTools; 

end PaveSet;
