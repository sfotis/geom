-- Created on: 2000-10-27
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CommonPrt from XIntTools 

	---Purpose: The class  is  to  describe a  common  part  
    	--          between two edges in  3-d space.

uses
    Edge  from  TopoDS, 
    ShapeEnum from  TopAbs, 
    Range  from  XIntTools,
    SequenceOfRanges  from  XIntTools, 
    Pnt from gp 
is 
    Create   
    	returns  CommonPrt from XIntTools; 
    	---Purpose: 
    	--- Empty constructor
    	---
     
    Create  (aCPrt:CommonPrt from XIntTools)   
    	returns  CommonPrt from XIntTools; 
    	---Purpose: 
    	--- Copy  constructor
    	---
     
    Assign  (me:out;  Other : CommonPrt from XIntTools) 
    	returns  CommonPrt from XIntTools;
    	---C++:  alias  operator = 
    	---C++:  return  & 
     
    SetEdge1  (me:out; anE:Edge from TopoDS); 	 
    	---Purpose:
    	--- Sets the first edge.
	---
    
    SetEdge2  (me:out; anE:Edge from TopoDS); 	 
    	---Purpose:  
    	--- Sets the second edge. 
	---
     
    SetType   (me:out; aType:ShapeEnum from  TopAbs); 
    	---Purpose:
    	--- Sets the type of  the common  part 
    	--- Vertex  or  Edge
	---

    SetRange1 (me:out;  aR: Range  from  XIntTools);
    	---Purpose: 
    	--- Sets the range of first edge. 
	---
     
    SetRange1 (me:out;  tf,tl: Real from Standard);
    	---Purpose: 
    	--- Sets the range of first edge.  
	---
     
    AppendRange2 (me:out;  aR: Range  from  XIntTools);
    	---Purpose: 
    	--- Appends the range of second edge.
	---
    
    AppendRange2 (me:out;  tf,tl: Real from Standard);
    	---Purpose: 
    	--- Appends the range of second edge.
	---
     
    SetVertexParameter1( me:out;  tV: Real from Standard);
    	---Purpose:
	--- Sets a parameter of first vertex
	---
     
    SetVertexParameter2( me:out;  tV: Real from Standard);
    	---Purpose:
	--- Sets a parameter of second vertex
	---

    Edge1     (me)   
    	returns Edge  from  TopoDS; 
    	---C++:  return  const& 
    	---Purpose: 
    	--- Returns the first edge.
	---
    
    Edge2     (me)   
    	returns Edge  from  TopoDS; 
    	---C++:  return  const&
    	---Purpose: 
    	--- Returns the second edge
	---
    
    Type      (me)   
    	returns  ShapeEnum from  TopAbs; 
    	---Purpose: 
    	--- Returns the type of  the common  part
	---
    
    Range1    (me)   
    	returns  Range  from  XIntTools;   
    	---C++:  return  const&
	---Purpose:
	--- Returns the range of first edge
	---
     
    Range1    (me; tf,tl:out Real from Standard);   
    	---Purpose: 
    	--- Returns the range of first edge. 
	---
     
    Ranges2   (me) 
    	returns  SequenceOfRanges from XIntTools; 
    	---C++:  return  const&  
    	---Purpose: 
    	--- Returns the  ranges of second edge.
	---
       
    ChangeRanges2   (me:out) 
    	returns  SequenceOfRanges from XIntTools; 
    	---C++:  return &  
    	---Purpose: 
    	--- Returns the  ranges of second edge.
	---
     
    VertexParameter1(me) 
    	returns Real from Standard;
	---Purpose:
	--- Returns parameter of first vertex
	---
      
    VertexParameter2(me) 
    	returns Real from Standard;
	---Purpose:
	--- Returns parameter of second vertex
	---
     
    Copy      (me;  anOther:out  CommonPrt from XIntTools); 
    	---Purpose: 
    	--- Copies me to anOther
	---
     
    AllNullFlag(me) 
        returns Boolean from Standard; 
	---Purpose:
	--- Modifier
	---
	 
    SetAllNullFlag(me:out; 
    	aFlag:Boolean from Standard); 
	---Purpose:
	--- Selector
	---

--
    SetBoundingPoints(me:out; 
	aP1: Pnt from gp;     
	aP2: Pnt from gp);
	---Purpose:
	--- Modifier
	---

    BoundingPoints(me; 
	aP1:out Pnt from gp;     
	aP2:out Pnt from gp);
	---Purpose:
	--- Selector
	---
--
fields
    myEdge1  :  Edge  from  TopoDS;
    myEdge2  :  Edge  from  TopoDS;
    myType   :  ShapeEnum from  TopAbs; 
    myRange1 :  Range  from  XIntTools;
    myVertPar1  :  Real from Standard;  
    myVertPar2  :  Real from Standard;  
    myRanges2:  SequenceOfRanges  from  XIntTools;

    myAllNullFlag: Boolean  from  Standard;
--
    myPnt1  :  Pnt from gp;
    myPnt2  :  Pnt from gp;
--

end CommonPrt;
