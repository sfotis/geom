-- Created on: 2002-02-04
-- Created by: Peter KURNEV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class WireShape from XBOP inherits Builder from XBOP

	---Purpose: 
    	--  The Root class to perform a Boolean Operations (BO)       
	--  Common,Cut,Fuse  between arguments when one of them is  
    	--  a wire          

uses
--    Wire   from TopoDS, 
    ListOfShape from TopTools

is 
    Create   
    	returns  WireShape from XBOP; 
    	---Purpose:  
    	--- Empty constructor;
    	---

    ---------------------------------------------- 
    --     
    --         W E S  C O M P O N E N T S  
    --     
    --            (for internal usage)    
    --     
    --      
    AddSplitPartsINOUT(me:out);   

    AddSplitPartsON(me:out);  

    MakeResult(me:out);   
    	---Purpose:   
    	--- Constructs the result of the BO 
    	---
     
    		    
fields 

    myLS        : ListOfShape from TopTools   
    	is protected;  

end WireShape;
