-- Created on: 2001-04-13
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class WESCorrector from XBOP 

	---Purpose: 
    	---  The algorithm to change the Wire Edges Set (WES) contents.
    	--   The NewWES will contain only wires instead of wires and edges. 
    	--
uses
    WireEdgeSet          from XBOP,
    PWireEdgeSet         from XBOP,
    ListOfConnexityBlock from XBOP 
    
is 
    Create   
    	returns WESCorrector from XBOP; 
    	---Purpose:  
    	--- Empty constructor; 
    	---
    SetWES  (me:out; 
		aWES: WireEdgeSet from XBOP);  
    	---Purpose: 
    	--- Modifier 
    	---
    Do (me:out); 
    	---Purpose: 
    	--- Performs the algorithm that  consists  of  two  steps 
    	--- 1. Make conexity blocks (  DoConnexityBlocks()  )     
    	--- 2. Make corrections     (  DoCorrections()  )        
    	---
    DoConnexityBlocks(me:out) 
    	is  private; 
       
    DoCorrections(me:out) 
    	is  private; 
      
    IsDone(me)  
    	returns Boolean from Standard;   
    	---Purpose: 
    	--- Selector 
    	---
    ErrorStatus	(me)  
    	returns Integer from Standard; 
    	---Purpose: 
    	--- Selector  
    	--- contents see XBOP_WESCorrector.cxx  
    	---
    WES     (me:out) 
    	returns WireEdgeSet from XBOP; 
    	---C++:  return &  
    	---Purpose: 
    	--- Selector 
    	---
    NewWES  (me:out) 
    	returns WireEdgeSet from XBOP; 
    	---C++:  return &   
    	---Purpose: 
    	--- Selector 
    	---

fields 

    myWES             : PWireEdgeSet         from XBOP; 
    myNewWES          : WireEdgeSet          from XBOP;  
    myConnexityBlocks : ListOfConnexityBlock from XBOP;  
    myIsDone          : Boolean from Standard;  
    myErrorStatus     : Integer from Standard;  

end WESCorrector;
