-- Created on: 2001-03-14
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CommonBlockAPI from XBOPTools 

	---Purpose:  
	--- class that provide some  useful tools 
    	--- to manage with a List Of Common Block-s             

uses
    ListOfCommonBlock from XBOPTools, 
    ListOfPaveBlock   from XBOPTools, 
    PaveBlock         from XBOPTools 
    
is 
    Create  (aList:ListOfCommonBlock from XBOPTools)   
    	returns CommonBlockAPI from XBOPTools; 
    	---Purpose:   
    	--- Constructor 
    	---
    List(me) 
    	returns  ListOfCommonBlock from XBOPTools; 
    	---C++:  return const & 
    	---Purpose:   
    	--- Selector 
    	---
    CommonPaveBlocks(me;   
    	    anE:Integer from  Standard) 
    	returns  ListOfPaveBlock from XBOPTools;
    	---C++:  return const &  
    	---Purpose:   
    	--- Returns all PaveBlock-s (from the list) that are 
    	--- common for the given edge with  DS-index <anE>     
    	---
    IsCommonBlock   (me;  
    	    aPB: PaveBlock from XBOPTools) 
    	returns  Boolean from Standard;
    	---Purpose:   
    	--- Returns TRUE if given PaveBlock <aPB> is 
    	--- common for the Blocks from the list      
    	---
fields 
    myListOfCommonBlock  :Address from Standard;
    myListOfPaveBlock    :ListOfPaveBlock from XBOPTools; 
    
end CommonBlockAPI;
