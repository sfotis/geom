-- Created on: 2001-05-28
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SolidStateFiller from XBOPTools  inherits StateFiller from XBOPTools 

	---Purpose:  
    	--  class to compute states (3D)  for the edges  (and theirs  
	--- split parts), vertices, wires, faces, shells  
        --- 
	 
	
uses 
    PPaveFiller from XBOPTools, 
    PaveFiller  from XBOPTools,  
    PShapesDataStructure from XBooleanOperations, 
    StateOfShape         from XBooleanOperations, 
    
    Shape from TopoDS,   
    Edge  from TopoDS, 
    
    State from TopAbs, 
     
    ShapeEnum from TopAbs
    
is 
    Create (aFiller: PaveFiller from XBOPTools) 
    	returns SolidStateFiller from XBOPTools; 
    	---Purpose:  
    	--- Constructor 
    	---
    Do(me:out)  
    	is redefined;
    	---Purpose: 
    	--- Launch the Filler   
    	---
    ---   
    --- 
    ---    private block 
    ---  
    DoNonSections  (me:out; 
    	    iRankShape: Integer from Standard) 
	is  private;  
    DoShellNonSections  (me:out; 
    	    iRankShape: Integer from Standard) 
	is  private; 

    DoSections  (me:out) 
	is  private; 

    IsFaceIntersected(me:out; 
    	    nF: Integer from Standard) 
    	returns Boolean from Standard 
    	is  private; 
     
end SolidStateFiller;
