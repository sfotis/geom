-- Created on: 2001-01-26
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class InterferencePool from XBOPTools 

	---Purpose:  
    	--  Class for storing information about  
    	--- results of all interferences for all shapes 

uses 
    ShapesDataStructure  from XBooleanOperations, 
    PShapesDataStructure from XBooleanOperations,  
    KindOfInterference   from XBooleanOperations, 
    
    CArray1OfInterferenceLine from XBOPTools, 
    CArray1OfSSInterference   from XBOPTools,
    CArray1OfESInterference   from XBOPTools,
    CArray1OfVSInterference   from XBOPTools, 
    CArray1OfEEInterference   from XBOPTools, 
    CArray1OfVEInterference   from XBOPTools, 
    CArray1OfVVInterference   from XBOPTools, 
    PShapeShapeInterference   from XBOPTools 
is 
    Create  
    	returns InterferencePool from XBOPTools ; 
    	---Purpose:  
    	--- Empty constructor 
    	---
    Create  (aDS:ShapesDataStructure from XBooleanOperations)
    	returns InterferencePool from XBOPTools ;  
    	---Purpose:   
    	--- Constructor 
    	---
    SetDS  (me:out;aDS:ShapesDataStructure from XBooleanOperations); 
    	---Purpose:  
    	--- Modifier  
    	---
    DS(me) 
    	returns  PShapesDataStructure from XBooleanOperations; 
    	---Purpose:  
    	--- Selector  
    	---
    HasInterference  (me; 
    	     anInd  :Integer from Standard) 
	returns Boolean from Standard;  
    	---Purpose: 
    	--- Returns  TRUE if the shape with DS_index  <anInd> 
    	--- has at least one  interference with non-empty result            
    	---
    IsComputed     (me;   
    	     anInd1  :  Integer from Standard;
    	     anInd2  :  Integer from Standard) 
	returns Boolean from Standard;  
    	---Purpose: 
    	--- Returns  TRUE if the interference between shapes  
    	--- <anInd1> and <anInd2> has already been computed.           
    	---
    SortTypes      (me;   
    	    	anInd1:in out Integer from Standard; 
                anInd2:in out Integer from Standard); 
    	---Purpose: 
    	--- Sorts types of shapes <anInd1> and <anInd2> in increasing order 
    	---
    InterferenceType  (me;   
    	    	anInd1: Integer from Standard; 
    	    	anInd2: Integer from Standard) 
    	returns KindOfInterference from XBooleanOperations;  
    	---Purpose: 
    	--- Gets the type of interference in accordance with the types of  
    	--- shapes  <anInd1> and <anInd2>
    	---
    AddInterference   (me:out;   
    	    	anInd1:  Integer from Standard;
    	    	anInd2:  Integer from Standard; 
                aType:   KindOfInterference from XBooleanOperations; 
	    	anIndex: Integer from Standard);  
    	---Purpose: 
    	--- Adds the info about interference in InterferenceLine-s for  
    	--- shapes  <anInd1> and <anInd2>
    	---
    InterferenceTable (me) 
    	returns  CArray1OfInterferenceLine from XBOPTools; 
    	---C++:  return  const& 
    	---Purpose: 
    	--- Returns the reference to complete array of interference line-s 
    	---
    SSInterferences (me:out)  
	returns CArray1OfSSInterference   from XBOPTools; 
    	---C++:  return  & 
    	---Purpose: 
    	--- Returns the reference to array Of F/F interferences 
    	---
    ESInterferences (me:out)  
	returns CArray1OfESInterference   from XBOPTools; 
    	---C++:  return  & 
    	---Purpose: 
    	--- Returns the reference to array Of E/F interferences 
    	---
    VSInterferences (me:out)  
	returns CArray1OfVSInterference   from XBOPTools; 
    	---C++:  return  &
    	---Purpose: 
    	--- Returns the reference to array Of V/F interferences 
    	---
    EEInterferences (me:out)  
	returns CArray1OfEEInterference   from XBOPTools; 
    	---C++:  return  &  
    	---Purpose: 
    	--- Returns the reference to arrray Of E/E interferences 
    	---
    VEInterferences (me:out)  
	returns CArray1OfVEInterference   from XBOPTools; 
    	---C++:  return  &  	 	
    	---Purpose: 
    	--- Returns the reference to arrray Of  V/E interferences 
    	---
    VVInterferences (me:out)  
	returns CArray1OfVVInterference   from XBOPTools; 
    	---C++:  return  &  	 	
    	---Purpose: 
    	--- Returns the reference to arrray Of  V/V interferences 
    	---
    -------------- 
    SSInterfs (me)  
	returns CArray1OfSSInterference   from XBOPTools; 
    	---C++:  return const & 
     
    ESInterfs (me)  
	returns CArray1OfESInterference   from XBOPTools; 
    	---C++:  return const & 
     
    VSInterfs (me)  
	returns CArray1OfVSInterference   from XBOPTools; 
    	---C++:  return const &
     
    EEInterfs (me)  
	returns CArray1OfEEInterference   from XBOPTools; 
    	---C++:  return const &  
	    
    VEInterfs (me)  
	returns CArray1OfVEInterference   from XBOPTools; 
    	---C++:  return const &  	 	
		 
    VVInterfs (me)  
	returns CArray1OfVVInterference   from XBOPTools; 
    	---C++:  return const & 
     

    GetInterference (me; 
    	    anIndex:  Integer from Standard; 
            aType  :  KindOfInterference from XBooleanOperations) 
	returns PShapeShapeInterference from XBOPTools; 


fields 
 
    myDS               :  PShapesDataStructure from XBooleanOperations;  
    myNbSourceShapes   :  Integer  from  Standard;  
    
    myInterferenceTable:  CArray1OfInterferenceLine from XBOPTools; 
    mySSInterferences  :  CArray1OfSSInterference   from XBOPTools;
    myESInterferences  :  CArray1OfESInterference   from XBOPTools;
    myVSInterferences  :  CArray1OfVSInterference   from XBOPTools;
    myEEInterferences  :  CArray1OfEEInterference   from XBOPTools;
    myVEInterferences  :  CArray1OfVEInterference   from XBOPTools;
    myVVInterferences  :  CArray1OfVVInterference   from XBOPTools;

end InterferencePool;
