-- Created on: 2001-04-09
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class EdgeInfo from XBOP 

    	---Purpose: 
    	---  The  auxiliary class to store data about edges 
    	---  that have common vertex         	 
	--- 
uses
    Edge from TopoDS 
    
--raises

is 
    Create 
    	returns EdgeInfo from XBOP;
    	---Purpose:  
    	--- Empty constructor;  
    	---
    SetEdge   (me:out; 
    	        aE:Edge from TopoDS); 
    	---Purpose: 
    	--- Modifier
    	---
    SetPassed (me:out;   
    	        aFlag:Boolean from Standard); 
    	---Purpose: 
    	--- Modifier
    	---
    SetAngle  (me:out;   
    	        anAngle:Real from Standard);  
    	---Purpose: 
    	--- Modifier
    	---
    SetInFlag (me:out;   
    	        aFlag:Boolean from Standard); 
    	---Purpose: 
    	--- Modifier
    	---
    Edge      (me) 
    	returns Edge from TopoDS; 
    	---C++:  return const & 
    	---Purpose: 
    	--- Selector
    	---
    Passed    (me) 
	returns Boolean from Standard; 
    	---Purpose: 
    	--- Selector
    	---
    Angle     (me) 
	returns Real from Standard;      
    	---Purpose: 
    	--- Selector
    	---
    IsIn      (me) 
    	returns Boolean from Standard;  
    	---Purpose: 
    	--- Selector
    	---
fields  

    myEdge  : Edge from TopoDS; 
    myPassed: Boolean from Standard; 
    myInFlag: Boolean from Standard; 
    myAngle : Real from Standard;     
     
end EdgeInfo;
