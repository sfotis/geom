-- Created on: 2000-11-21
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Interference from XBOPTools 

	---Purpose: class for storing information about an interference 
	---         that  takes  place  between  given  shape and shape 
        ---         with  DS-index =aWith  	 


uses
    KindOfInterference from XBooleanOperations

is 
    Create 
    	returns Interference from XBOPTools;  
    	---Purpose:  
    	--- Empty constructor 
    	---
    Create  (aWith   :Integer from Standard; 
    	     aType   :KindOfInterference from XBooleanOperations; 
	     anIndex :Integer from Standard)
    	returns Interference from XBOPTools;   
    	---Purpose:  constructor 
    	--- aWith  -  DS-index for the opposite shape     
    	--- aType  -  the type of the  interference       
    	--- anIndex-  the index of the result in corresponding  
    	--- interference table  (if the result is computed 
    	--- but there is no result  ->   anIndex=0) 
    	---
    SetWith  (me:out; aWith :Integer from Standard);	
    	---Purpose:  
    	--- Modifier 
    	---
    SetType  (me:out; aType : KindOfInterference from XBooleanOperations); 
    	---Purpose: 
    	--- Modifier 
    	---
    SetIndex (me:out; anIndex  :Integer from Standard); 
    	---Purpose: 
    	--- Modifier 
    	---
    With  (me) 
    	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector  
    	---
    Type  (me)  
    	returns  KindOfInterference from XBooleanOperations; 
    	---Purpose:  
    	--- Selector  
    	---
    Index (me) 
    	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector  
    	---

fields
    myWith        : Integer from Standard; 
    myType        : KindOfInterference from XBooleanOperations; 
    myIndex       : Integer from Standard;  --< index  in corresp.interference  table  
   

end Interference;
