-- Created on: 2001-12-24
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Refiner from XBOP 

	---Purpose:  
	--  The  algorithm to provide the refinition  
    	--  for a resulting shape of Boolean Operation  
    	--  algorithm.   
        --  (not  completed  yet)	     


uses
    Shape from TopoDS,
    ListOfShape from TopTools 
    
--raises

is 
    Create   
    	returns Refiner from XBOP; 
    	---Purpose:  
    	--- Empty constructor;  
    	---
    Create(aS: Shape from TopoDS)    
    	returns Refiner from XBOP; 
    	---Purpose:  
    	--- Constructor;  
    	---
    SetShape(me:out; 
    	   aS: Shape from TopoDS); 
    	---Purpose: 
    	--- Modifier
    	---
    SetInternals (me:out; 
	   aLS:ListOfShape from TopTools); 
    	---Purpose: 
    	--- Modifier
    	---
    Do(me:out); 
    	---Purpose: 
    	--- Performs the algorithm  
    	---
    IsDone(me) 
    	returns Boolean from Standard; 
    	---Purpose: 
    	--- Selector
    	---
    ErrorStatus(me) 
    	returns Integer from Standard; 
    	---Purpose: 
    	--- Selector
    	---
    Shape(me) 
    	returns Shape from TopoDS; 
    	---C++: return const & 
    	---Purpose: 
    	--- Selector
    	---
    NbRemovedVertices(me) 
 	 returns Integer from Standard; 
    	---Purpose: 
    	--- Selector
    	---
    NbRemovedEdges(me) 
 	 returns Integer from Standard;  
    	---Purpose: 
    	--- Selector
    	---
    DoInternals(me:out) is  private; 
    	---Purpose: 
    	--- Internal usage
    	---


fields
 
    myShape       : Shape   from TopoDS; 
    myIsDone      : Boolean from Standard; 
    myErrorStatus : Integer from Standard;	     
    myNbRemovedVertices  : Integer from Standard;	
    myNbRemovedEdges     : Integer from Standard;	 
    myInternals   : ListOfShape from TopTools; 
    
end Refiner;
