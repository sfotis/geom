-- Created on: 2005-10-05
-- Created by: Mikhail KLOKOV
-- Copyright (c) 2005-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class CurveRangeSample from XIntTools inherits BaseRangeSample from XIntTools
uses
    Range from XIntTools
is

    Create
    	returns CurveRangeSample from XIntTools;

    Create(theIndex: Integer from Standard)
    	returns CurveRangeSample from XIntTools;

    SetRangeIndex(me: in out; theIndex: Integer from Standard);
	---C++: inline

    GetRangeIndex(me)
    	returns Integer from Standard;
	---C++: inline
	
    IsEqual(me; Other: CurveRangeSample from XIntTools)
    	returns Boolean from Standard;
	---C++: inline

    GetRange(me; theFirst, theLast: Real from Standard; 
    	    	 theNbSample: Integer from Standard)
    	returns Range from XIntTools;

    GetRangeIndexDeeper(me; theNbSample: Integer from Standard)
    	returns Integer from Standard;
	---C++: inline

fields
    myIndex: Integer from Standard;

end CurveRangeSample from XIntTools;
