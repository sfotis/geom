-- Created on: 2001-02-15
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PaveBlock from XBOPTools 

	---Purpose:  
    	--  Class for storing info about a couple  
        --- of neighbouring paves on an edge  

uses
    Pave from XBOPTools,  
    PointBetween from XBOPTools,
    Range        from XIntTools, 
    ShrunkRange  from XIntTools, 
    Curve        from XIntTools



is 
    Create 
    	returns PaveBlock from XBOPTools;  
    	---Purpose: 
    	--- Empty constructor 
    	---
    Create (anEdge:  Integer from Standard; 
    	    aPave1:  Pave from XBOPTools; 
    	    aPave2:  Pave from XBOPTools); 
    	---Purpose:  
    	--- Constructor 
    	--- Index  - DS-index of the edge    	 
    	--- aPave1 - one pave              
    	--- aPave2 - other pave               
    	---
    SetEdge (me:out;   
    	     anEdge:Integer from Standard); 
    	---Purpose:  
    	--- Modifier  
    	--- Sets DS-index for the edge that is between aPave1 and aPave2 
    	---
    SetOriginalEdge  (me:out;   
    	    	      anEdge:Integer from Standard);  
    	---Purpose:  
    	--- Modifier  
    	--- Sets DS-index for the edge from which this pave block comes from 
    	---
    SetPave1(me:out;  
    	     aPave: Pave from XBOPTools);	     
    	---Purpose:  
    	--- Modifier  
    	---
    SetPave2(me:out;  
    	     aPave: Pave from XBOPTools);	     
    	---Purpose:  
    	--- Modifier  
    	---
    SetShrunkRange  (me:out;   
    	    	     aSR:ShrunkRange from XIntTools);  
    	---Purpose:  
    	--- Modifier  
    	--- Sets the Shrunk Range for the pave block 
    	---
    SetPointBetween (me:out; 
    	    	     aP: PointBetween from XBOPTools);  
    	---Purpose:  
    	--- Modifier  
    	--- Sets the point between the paves for the pave block  
    	---

    ---  Case  of  Face/Face Pave  Block 
    ---		    	     
    SetCurve        (me:out; 
    	    	     aC:Curve from XIntTools);  
    	---Purpose:  
    	--- Modifier  
    	--- Sets the intersection curve to which the pave block belongs to  
    	---
    SetFace1        (me:out; 
    	    	     nF1:Integer from Standard); 
    	---Purpose:  
    	--- Modifier  
    	--- Sets the DS-index of the first face  
    	---
    SetFace2        (me:out; 
    	    	     nF2:Integer from Standard);  
    	---Purpose:  
    	--- Modifier  
    	--- Sets the DS-index of the second face  
    	---
    Edge    (me) 
    	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector  
    	---
    OriginalEdge(me) 
    	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector  
    	---
    Pave1(me) 
    	returns Pave from XBOPTools; 
    	---C++:  return const &	 
    	---Purpose:  
    	--- Selector  
    	---
    Pave2(me) 
    	returns Pave from XBOPTools; 
    	---C++:  return const &	
    	---Purpose:  
    	--- Selector  
    	---
    IsValid(me) 
	returns Boolean from Standard;	    	     
    	---Purpose:  
    	--- Returns  TRUE if both paves have vertex index !=0            
    	---
    IsEqual(me;  
    	    Other:PaveBlock from XBOPTools)    
        returns Boolean from Standard;	
    	---Purpose:  
    	--- Returns  TRUE if <Other> is  equal to me 
    	---
    Parameters   (me; 
                  aT1:out Real from Standard;   
                  aT2:out Real from Standard);    
    	---Purpose:  
    	--- Returns values for paves' parameters      
    	---
    Range  (me) 
    	returns Range from XIntTools; 
    	---C++:  return const &	
    	---Purpose:  
    	--- Returns parmetric range for paves' parameters      
    	---
    ShrunkRange(me) 
    	returns ShrunkRange from XIntTools; 
    	---C++:  return const &  
    	---Purpose:  
    	--- Selector      
    	---
    PointBetween  (me) 
    	returns  PointBetween from XBOPTools; 
    	---C++:  return const & 	 
    	---Purpose:  
    	--- Selector      
    	---
    Curve(me) 
    	returns Curve from XIntTools; 
    	---C++:  return const & 
    	---Purpose:  
    	--- Selector      
    	---
    Face1(me) 
    	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector      
    	---
    Face2(me) 
    	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector      
    	---
    IsInBlock(me; 
    	   aPaveX:  Pave from XBOPTools) 
    	returns Boolean  from Standard;  
    
fields   

    myEdge         :  Integer from Standard;
    myOriginalEdge :  Integer from Standard;
    myPave1        :  Pave from XBOPTools; 
    myPave2        :  Pave from XBOPTools; 
    myRange        :  Range from XIntTools;     
    myShrunkRange  :  ShrunkRange from XIntTools; 
    myCurve        :  Curve from XIntTools; 
    myFace1        :  Integer from Standard; 
    myFace2        :  Integer from Standard; 
    myPointBetween :  PointBetween from XBOPTools;  
     
end PaveBlock;
