-- Created on: 2001-04-17
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class CorrectTolerances from XBOP 

    	---Purpose: 
	---  The  Set  of  static functions to provide valid values of  
    	---  tolerances for shapes.     
    	---  Tolerances becomes valid in  terms of the checkshape.    

uses
    Shape  from  TopoDS 
    
is 
    CorrectTolerances      (myclass;  
    	    	    	    aS: Shape  from  TopoDS; 
    	    	    	    aTolMax: Real from Standard =0.0001);  
    	---Purpose:	 
    	--- Provides valid values of tolerances for the shape <aS>         
    	--- <aTolMax> is max value of the tolerance that can be 
    	--- accepted for correction.  If real value of the tolerance 
    	--- will be greater than  <aTolMax>, the correction does not 
    	--- perform. 
    	---
    CorrectCurveOnSurface  (myclass;  
    	    	    	    aS: Shape  from  TopoDS; 
    	    	    	    aTolMax: Real from Standard =0.0001); 
    	---Purpose:	 
    	--- Provides valid values of tolerances for the shape <aS> 
    	--- in  terms of BRepCheck_InvalidCurveOnSurface.   
    	---
    CorrectPointOnCurve    (myclass;  
    	    	    	    aS: Shape  from  TopoDS; 
    	    	    	    aTolMax: Real from Standard =0.0001);  		    
    	---Purpose:	 
    	--- Provides valid values of tolerances for the shape <aS> 
    	--- in  terms of BRepCheck_InvalidPointOnCurve.   
    	---

end CorrectTolerances;
