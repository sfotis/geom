-- Created on: 2004-09-02
-- Created by: Oleg FEDYAEV
-- Copyright (c) 2004-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class CheckResult from XBOPTools
    ---Purpose: contains information about faulty shapes
    --          and faulty types
uses 
    
    Shape       from TopoDS,
    ListOfShape from TopTools,
    CheckStatus from XBOPTools,
    Geometry    from Geom

is

    Create
    	returns CheckResult;
    ---Purpose: empty constructor

    AddShape(me: in out; TheShape: Shape from TopoDS);
    ---Purpose: adds a shape with faulty to a list

    GetShapes(me)
    	returns ListOfShape from TopTools;
    ---C++: return const &
    ---Purpose: gets access to faulty shapes in a list const

    SetCheckStatus(me:in out; TheStatus: CheckStatus from XBOPTools);
    ---Purpose: sets faulty status for shapes

    GetCheckStatus(me)
    	returns  CheckStatus from XBOPTools;
    ---Purpose: gets faulty status for shapes

    SetInterferenceGeometry(me: in out; TheGeometry: Geometry from Geom);
    ---Purpose: sets an attached geometry to faulty shapes if any

    GetInterferenceGeometry(me)
    	returns Geometry from Geom;
    ---C++: return const &
    ---Purpose: gets an attached geometry to shapes if any

fields

    myStatus   : CheckStatus from XBOPTools;
    myShapes   : ListOfShape from TopTools;
    myGeometry : Geometry    from Geom;

end CheckResult;
