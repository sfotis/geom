-- Created on: 1995-12-21
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

--modified by NIZNHY-PKV Tue Apr  3 15:53:58 2001   

class FaceAreaBuilder from XBOP inherits Area2dBuilder from XBOP

    ---Purpose: 
    -- The FaceAreaBuilder algorithm is used to construct Faces from a LoopSet,
    -- where the Loop is the composite topological object of the boundary,
    -- here wire or block of edges.
    -- The LoopSet gives an iteration on Loops.
    -- For each Loop  it indicates if it is on the boundary (wire) or if it
    -- results from  an interference (block of edges).
    -- The result of the FaceAreaBuilder is an iteration on areas.
    -- An area is described by a set of Loops.

uses

    LoopSet        from XBOP,
    LoopClassifier from XBOP
    
is

    Create returns FaceAreaBuilder;
    	---Purpose:  
    	--- Empty constructor; 
    	---
    Create(LS :out LoopSet from XBOP;  
    	   LC :out LoopClassifier from XBOP;
    	   ForceClass : Boolean = Standard_False)  
    	returns FaceAreaBuilder;
    	---Purpose:  
    	--- Creates the object to build faces on the (wires,blocks of edge)  
    	--- of <LS>, using the classifier <LC>.
	---
    InitFaceAreaBuilder(me :out;
    	    	   	LS :out LoopSet from XBOP;  
    	    	        LC :out LoopClassifier from XBOP;
    	    	    	ForceClass : Boolean = Standard_False) 
    	 is static;
    	---Purpose:  
    	--- Initializes the object to build faces on the (wires,blocks of edge)  
    	--- of <LS>, using the classifier <LC>.
	---
end FaceAreaBuilder;
