-- Created on: 2000-11-21
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class VSInterference from XBOPTools 
    inherits ShapeShapeInterference from XBOPTools  
    
    	---Purpose:  
    	--  Class for storing info about an Verex/Face interference
	--- 
is
    Create  
    	returns  VSInterference from XBOPTools; 
    	---Purpose:  
    	--- Empty constructor  
    	---
    Create  (anIndex1:  Integer from Standard;  
    	     anIndex2:  Integer from Standard; 
    	     U: Real from Standard;  
    	     V: Real from Standard)
    	returns  VSInterference from XBOPTools;  
    	---Purpose:   
    	--- Constructor  
    	--- anIndex1,  
    	--- anIndex2 see XBOPTools_ShapeShapeInterference for details      
    	--- U, V  -  values of parameters on the surface    
    	---
    SetUV   (me:out; U, V: Real from Standard); 
    	---Purpose:  
    	--- Modifier   
    	---
    UV      (me;  U:out Real from Standard;   
                  V:out Real from Standard);
    	---Purpose:  
    	--- Selector  
    	---
fields
    myU:Real from Standard;  
    myV:Real from Standard;  

end VSInterference;
