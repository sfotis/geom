-- Created on: 1995-12-21
-- Created by: Jean Yves LEBEY 
-- Copyright (c) 1995-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.

-- modified by PKV Tue Apr  3 16:57:39 2001


class FaceBuilder from XBOP 

    ---Purpose: 
    ---   The  algorithm to   construct Faces from a WireEdgeSet        
    --- 
    
uses

    Shape  from TopoDS,
    Face   from TopoDS, 
    Wire   from TopoDS, 
    Edge   from TopoDS, 
    Vertex from TopoDS, 
    ListOfShape from TopTools, 
    SequenceOfInteger from TColStd,  
    Context from XIntTools,
    WireEdgeSet     from XBOP,
    PWireEdgeSet    from XBOP
--    LoopSet         from XBOP,
--    BlockIterator   from XBOP,
--    BlockBuilder    from XBOP,
--    FaceAreaBuilder from XBOP, 
   

is

    Create  
    	returns FaceBuilder;
    	---Purpose:  
    	--- Empty constructor; 
    	---
    Do(me :out;  
    	   aWES        : WireEdgeSet from XBOP;  
    	   aForceClass : Boolean from Standard =Standard_True); 
    	---Purpose: 
    	--- Launches the algorithm consisting of four steps 
    	--- 1.  Split the WES on wires       
    	--- 2.  Make Loops from wires         
    	--- 3.  Make Areas from Loops           
    	--- 4.  Make Faces from Areas    
    	---
    
    	---
--    BuildNewFaces (me :out) 
--    	is private;  
    	---Purpose:     
    	--- Make Faces from Areas  
    	--- 
 
--modified by NIZNHY-PKV Wed Feb 29 10:57:40 2012f    
    SetContext(me:out; 
    	    aCtx:Context from XIntTools); 
	---Purpose:  
        -- Sets intersection context <aCtx>
	  
    Context(me) 
    	returns Context from XIntTools; 
    	---C++: return const & 
     	---Purpose:  
        -- Returns intersection context 
--modified by NIZNHY-PKV Wed Feb 29 10:57:52 2012t 
 
    WES (me) 
    	returns  WireEdgeSet from XBOP; 
    	---C++: return const &
    	---Purpose:     
    	--- Selector 
    	---
    NewFaces (me) 
	returns ListOfShape from TopTools; 
    	---C++: return const &	
    	---Purpose:     
    	--- Selector 
    	---
    SetTreatment (me: out; 
	aTreatment: Integer from Standard);  
    	---Purpose:     
    	--- Modifier 
    	--- 0 -Treat internal edges,  
    	--- 1 -Do not treat internal edges      
    	---

    SetTreatSDScales (me: out; 
	aTreatment: Integer from Standard);  
    	---Purpose:     
    	--- Modifier 
    	--- 1 -Treat scale configured same domain faces,  
    	--- 0 -Do not treat them.     
	--- 
--    SetManifoldFlag(me: out; 
--    	aMFlag:  Boolean from Standard); 
    	---Purpose:     
    	--- Modifier 
    	---  
--    ManifoldFlag(me) 
--    	returns Boolean from Standard; 
    	---Purpose:     
    	--- Selector 
    	---
    Treatment (me) 
	returns Integer from Standard; 
    	---Purpose:     
    	--- Selector 
    	---
    TreatSDScales (me) 
	returns Integer from Standard; 
    	---Purpose:     
    	--- Selector 
    	---
    --- 
    --- 
    --- Faces' iterator   
    --- 
--    InitFace(me:out)  
--    	returns Integer from Standard;
    
--    MoreFace(me)  
--    	returns Boolean from Standard;
    
--    NextFace(me:out);
    ---Purpose:     
    --- 
    --- 
    --- Wires' iterator 
    ---  
--    InitWire(me:out)  
--    	returns Integer from Standard;
     
--    MoreWire(me)  
--    	returns Boolean from Standard;
     
--    NextWire(me:out); 
    	
--    IsOldWire(me)  
--    	returns Boolean from Standard;
     
--    OldWire(me)  
--    	returns Shape from TopoDS;
 --   	---C++: return const &
   
--    Wire(me)  
--    	returns Wire from TopoDS;
--    	---C++: return const &
--    	---Purpose:      
--    	---  

    ---  
    ---  Edges' iterator 
    ---
--    FindNextValidElement(me:out);
         
--    InitEdge(me:out)  
--    	returns Integer from Standard;
     
--    MoreEdge(me)  
--    	returns Boolean from Standard;
     
--    NextEdge(me : in out);
     
--    Edge(me)  
--    	returns Edge from TopoDS;
--    	---C++: return const &
    	---Purpose:      
    	--- 
	
--    MakeLoops(me :out; 
--    	      SS :out WireEdgeSet from XBOP) 
--    	is protected;
    	---Purpose:      
    	--- Make Loops from wires     
    	---
   DoInternalEdges (me :out) 
    	is protected;       		    	    
    	---Purpose:  
    	--- Processes internal edges if they exists     
    
    SDScales(me :out) 
    	is  protected; 
    	---Purpose:   
    	--- Treatment SD faces with a "scale" 
    	---
    --modified by NIZNHY-PKV Wed Feb 29 09:12:17 2012f 
    PerformAreas(me :out; 
    	      SS :out WireEdgeSet from XBOP) 
    	is protected; 
    --modified by NIZNHY-PKV Wed Feb 29 09:12:20 2012t 
    
fields

    myFace             : Face from TopoDS;
--    myLoopSet          : LoopSet         from XBOP;
--    myBlockIterator    : BlockIterator   from XBOP;
--    myBlockBuilder     : BlockBuilder    from XBOP;
--    myFaceAreaBuilder  : FaceAreaBuilder from XBOP;
    myWES              : PWireEdgeSet    from XBOP;
    myNewFaces         : ListOfShape     from TopTools; 
    myTreatment        : Integer from Standard;           
--    myManifoldFlag     : Boolean from Standard;     
    myTreatSDScales    : Integer from Standard;   
    myNegatives        : SequenceOfInteger from TColStd; 
    myContext          : Context from XIntTools; 
end FaceBuilder;
