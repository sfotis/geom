-- Copyright (C) 2007-2013  CEA/DEN, EDF R&D, OPEN CASCADE
--
-- Copyright (C) 2003-2007  OPEN CASCADE, EADS/CCR, LIP6, CEA/DEN,
-- CEDRAT, EDF R&D, LEG, PRINCIPIA R&D, BUREAU VERITAS
--
-- This library is free software; you can redistribute it and/or
-- modify it under the terms of the GNU Lesser General Public
-- License as published by the Free Software Foundation; either
-- version 2.1 of the License.
--
-- This library is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the GNU
-- Lesser General Public License for more details.
--
-- You should have received a copy of the GNU Lesser General Public
-- License along with this library; if not, write to the Free Software
-- Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301  USA
--
-- See http://www.salome-platform.org/ or email : webmaster.salome@opencascade.com
--

-- File:	NMTTools.cdl
-- Created:	Thu Dec  4 16:55:49 2003
-- Author:	Peter KURNEV
--		<pkv@irinox>
--
package NMTTools

	---Purpose:

uses

    TCollection,
    TColStd,
    gp,
    TopAbs,
    TopoDS,
    TopTools,
    Geom2d,
    XBooleanOperations,
    XBOPTColStd,
    XIntTools,
    XBOPTools,
    NMTDS

is
    imported CoupleOfShape from NMTTools;
    imported CommonBlock from NMTTools;
    imported CommonBlockAPI from NMTTools;
    imported FaceInfo from NMTTools;
    imported Tools from NMTTools;
    imported PaveFiller from NMTTools;
    imported PPaveFiller from NMTTools;
    imported DEProcessor from NMTTools;
    imported CheckerSI from NMTTools;
    --
    imported ListOfCommonBlock from NMTTools;
    imported ListIteratorOfListOfCommonBlock from NMTTools;

    imported ListOfCoupleOfShape from NMTTools;
    imported ListIteratorOfListOfCoupleOfShape from NMTTools;

    imported MapOfPaveBlock from NMTTools;
    imported MapIteratorOfMapOfPaveBlock from NMTTools;

    imported IndexedDataMapOfIndexedMapOfInteger from NMTTools;
    imported IndexedDataMapOfShapePaveBlock from NMTTools;
    imported IndexedDataMapOfShapeIndexedMapOfShape from NMTTools;

    imported DataMapOfIntegerListOfPaveBlock from NMTTools;
    imported DataMapIteratorOfDataMapOfIntegerListOfPaveBlock from NMTTools;

    imported DataMapOfIntegerFaceInfo from NMTTools;
    imported DataMapIteratorOfDataMapOfIntegerFaceInfo from NMTTools;

    imported CommonBlockPool from NMTTools;

    --
    --class PaveFiller;
    --class Tools;
    --class CommonBlock;
    --class CommonBlockAPI;
    --class FaceInfo;
    --class CoupleOfShape;
    --class CheckerSI;
    --class DEProcessor;
    --pointer PPaveFiller to PaveFiller from NMTTools;
    --
    --class ListOfCommonBlock  instantiates
    --	List from TCollection(CommonBlock from NMTTools);

    --class ListOfCoupleOfShape  instantiates
    --	List from TCollection(CoupleOfShape from NMTTools);
--
    --class  MapOfPaveBlock  instantiates
    --	Map from TCollection   (PaveBlock from XBOPTools,
    --	    	    	    	PaveBlockMapHasher from XBOPTools);
--
    --class IndexedDataMapOfIndexedMapOfInteger instantiates
    --	IndexedDataMap from TCollection  (Integer from Standard,
    --	    	    	    	    	  IndexedMapOfInteger from TColStd,
    --	    	    	    	    	  MapIntegerHasher from TColStd);

    --class IndexedDataMapOfShapePaveBlock instantiates
    --	IndexedDataMap from TCollection  (Shape from TopoDS,
    --	    	    	    	    	  PaveBlock from XBOPTools,
    --	    	    	    	    	  ShapeMapHasher from TopTools);

    --class IndexedDataMapOfShapeIndexedMapOfShape instantiates
    --	IndexedDataMap from TCollection  (Shape from TopoDS,
    --	    	    	    	    	  IndexedMapOfShape from TopTools,
    --	    	    	    	    	  ShapeMapHasher from TopTools);

--
    --class DataMapOfIntegerListOfPaveBlock instantiates
    --	DataMap from TCollection(Integer from  Standard,
    --	    	    	    	 ListOfPaveBlock from XBOPTools,
    --				 MapIntegerHasher from TColStd);

    --class DataMapOfIntegerFaceInfo instantiates
    --	DataMap from TCollection(Integer from  Standard,
    --                             FaceInfo from  NMTTools,
    --				 MapIntegerHasher from TColStd);
--
    --class CommonBlockPool    instantiates
    --	CArray1 from XBOPTColStd (ListOfCommonBlock from NMTTools);
--
end NMTTools;
