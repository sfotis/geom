-- Created on: 2001-09-12
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DEInfo from XBOPTools 

	---Purpose:  
    	--  Auxiliary class for storing  information about  
    	--- a degenerated edge 
      	---  

uses 
    ListOfInteger from TColStd

is 
    Create 
    	returns DEInfo from XBOPTools;
    	---Purpose:  
    	--- Empty constructor 
    	---
    SetVertex   (me:out; 
    	    nV:Integer from Standard); 
    	---Purpose: 
    	--- Modifier
    	--- Sets  DS-index for the vertex to which 
    	--- degenerated edge belongs to 	      
    	---
    SetFaces  	(me:out; 
    	    aLF: ListOfInteger from TColStd); 
    	---Purpose:  
    	--- Modifier
    	--- Sets  DS-indices for the faces to which 
    	--- degenerated edge belongs to    
    	---
    Faces(me) 
    	returns ListOfInteger from TColStd; 
    	---C++:  return const & 
    	---Purpose:  
    	--- Selector
    	---
    ChangeFaces(me:out) 
    	returns ListOfInteger from TColStd; 
    	---C++:  return & 
    	---Purpose:  
    	--- Selector/Modifier
    	---
    Vertex(me) 
    	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector
    	---

fields 
    myFaces  :  ListOfInteger from TColStd; 
    myVertex :  Integer from Standard; 
     
end DEInfo;
