-- Created on: 2001-06-25
-- Created by: Michael KLOKOV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class SolidAreaBuilder from XBOP inherits Area3dBuilder from XBOP

    	---Purpose: 
    	---   construct Areas for Solids from a Shell Faces Set        
	---
uses
    LoopSet        from XBOP,
    LoopClassifier from XBOP

is
    Create returns SolidAreaBuilder from XBOP;
    	---Purpose:  
    	--- Empty constructor; 
    	---
    Create(LS:out LoopSet from XBOP;
    	   LC:out LoopClassifier from XBOP;
	   ForceClassFlag: Boolean from Standard = Standard_False)
    	returns SolidAreaBuilder from XBOP;
    	---Purpose:  
    	--- Creates an  object to build solids on
    	--- the (shells,  blocks of faces) of <LS>,  
    	--- using the classifier <LC>.  
    
    InitSolidAreaBuilder(me: in out; 
    	    	    LS:out LoopSet from XBOP;
    	    	    LC:out LoopClassifier from XBOP;
		    ForceClassFlag: Boolean from Standard); 
    	---Purpose:   
    	---Purpose:  
    	--- Initialize the object to find the areas of
    	--- the shapes described by <LS>, 
    	--- using the classifier <LC>.   
    	---
end SolidAreaBuilder from XBOP;
