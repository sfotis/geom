-- Created on: 2001-09-12
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class DEProcessor from XBOPTools 

	---Purpose:  
    	--   
    	--  The  Algorithm to compute and store in interferences' pool 
	--- and in the Data  Structure  the following values        
    	--- for degenerated edges 
	---         1.  Paves/Pave set(s)
	---         2.  Split parts 
	---         3.  States (3D) for split parts 
        --- 
	
uses  

    Vertex from TopoDS,
    Edge   from TopoDS, 
    Face   from TopoDS, 
     
    PPaveFiller     from XBOPTools, 
    PaveFiller      from XBOPTools,   
    ListOfPaveBlock from XBOPTools,
     
    PShapesDataStructure from XBooleanOperations, 
    
    IndexedDataMapOfIntegerDEInfo from XBOPTools	  



is
    Create (aFiller: PaveFiller from XBOPTools; 
    	    aDim  : Integer from Standard=3) 
    	returns  DEProcessor from XBOPTools; 
    	---Purpose:  
    	--- Constructor 
    	---
    Do(me:out);   
    	---Purpose: 
    	--- Launches the processor   
    	---
    IsDone(me) 
    	returns Boolean from Standard; 
    	---Purpose:  
    	--- Returns TRUE if it is Ok       
    	---
    --- 
    ---    Private block 
    ---
    ---
    FindDegeneratedEdges (me:out) 
    	is  private; 
	
    DoPaves  (me:out) 
    	is  private; 
	 
    FindPaveBlocks (me:out; 
    	    nED:Integer from Standard; 
    	    nVD:Integer from Standard; 
    	    nFD:Integer from Standard; 
    	    aLPB:out ListOfPaveBlock from XBOPTools) 
    	is  private; 
     
    FillPaveSet (me:out; 
    	    nED:Integer from Standard; 
    	    nVD:Integer from Standard; 
    	    nFD:Integer from Standard; 
    	    aLPB:out ListOfPaveBlock from XBOPTools) 
    	is  private; 

    FillSplitEdgesPool(me:out; 
    	    nED:Integer from Standard)
    	is  private; 
  
    MakeSplitEdges(me:out; 
    	    nED:Integer from Standard;
    	    nFD:Integer from Standard)
    	is  private;   
	 
    MakeSplitEdge  (me:out;   
        	    aS1: Edge from TopoDS; 
		    aF : Face from TopoDS;	     
		    aV1: Vertex from TopoDS;	     
   	    	    aP1: Real from Standard; 
    	    	    aV2: Vertex from TopoDS; 
		    aP2: Real from Standard; 
    	    	    aNewEdge:out Edge from TopoDS) 
    	is  private; 		
     
    DoStates  (me:out; 
    	    nED:Integer from Standard;
    	    nFD:Integer from Standard)
    	is  private;    
	 
    DoStates2D  (me:out; 
    	    nED:Integer from Standard;
    	    nFD:Integer from Standard)
    	is  private; 
	 
fields 
    myDim     : Integer from Standard;     
    
    myFiller  : PPaveFiller from XBOPTools; 
    myDS      : PShapesDataStructure from XBooleanOperations;
    myIsDone  : Boolean   from Standard;   
    myDEMap   : IndexedDataMapOfIntegerDEInfo from XBOPTools; 
       
	     
end DEProcessor;
