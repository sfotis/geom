-- Created on: 2001-07-06
-- Created by: Michael KLOKOV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class BeanBeanIntersector from XIntTools

    ---Purpose: The class BeanBeanIntersector computes ranges of parameters on
    ---         the curve of a first bean (part of edge) that bounds the parts of bean which
    ---	        are on the other bean according to tolerance of edges.

uses
    SequenceOfRoots     from XIntTools,
    MarkedRangeSet      from XIntTools,
    SequenceOfRanges    from XIntTools,
    Range               from XIntTools,
    ExtCC               from Extrema,
    ProjectPointOnCurve from GeomAPI,
    Edge                from TopoDS,
    Curve               from BRepAdaptor,
    Curve               from Geom


is
    Create returns BeanBeanIntersector from XIntTools;
    
    Create(theEdge1: Edge from TopoDS;
    	   theEdge2: Edge from TopoDS)
	   returns BeanBeanIntersector from XIntTools;
    	---Purpose: 
    	--- Initializes the algorithm
	---

    Create(theCurve1        : Curve   from BRepAdaptor;
    	   theCurve2        : Curve from BRepAdaptor;
    	   theBeanTolerance1: Real from Standard;
    	   theBeanTolerance2: Real from Standard)
	   returns BeanBeanIntersector from XIntTools;
    	---Purpose: 
    	--- Initializes the algorithm
	---

    Create(theCurve1          : Curve   from BRepAdaptor;
    	   theCurve2          : Curve   from BRepAdaptor;
	   theFirstParOnCurve1: Real from Standard;
	   theLastParOnCurve1 : Real from Standard;
    	   theFirstParOnCurve2: Real from Standard;
	   theLastParOnCurve2 : Real from Standard;
    	   theBeanTolerance1  : Real from Standard;
    	   theBeanTolerance2  : Real from Standard)
	   returns BeanBeanIntersector from XIntTools;
    	---Purpose: 
    	--- Initializes the algorithm
	---

    Init(me: in out;theEdge1: Edge from TopoDS;
    	            theEdge2: Edge from TopoDS);
    	---Purpose: 
    	--- Initializes the algorithm
	---



    Init(me: in out;theCurve1        : Curve   from BRepAdaptor;
	    	    theCurve2        : Curve from BRepAdaptor;
    	    	    theBeanTolerance1: Real from Standard;
    	    	    theBeanTolerance2: Real from Standard);
    	---Purpose: 
    	--- Initializes the algorithm
	---

    Init(me: in out;theCurve1          : Curve   from BRepAdaptor;
    	    	    theCurve2          : Curve   from BRepAdaptor;
	    	    theFirstParOnCurve1: Real from Standard;
	    	    theLastParOnCurve1 : Real from Standard;
    	    	    theFirstParOnCurve2: Real from Standard;
	    	    theLastParOnCurve2 : Real from Standard;
    	    	    theBeanTolerance1  : Real from Standard;
    	    	    theBeanTolerance2  : Real from Standard);
    	---Purpose: 
    	--- Initializes the algorithm
	---

    SetBeanParameters(me: in out;IsFirstBean       : Boolean from Standard;
    	    	    	    	 theFirstParOnCurve: Real from Standard;
	    	    	    	 theLastParOnCurve : Real from Standard);
    	---Purpose: 
    	--- Sets bounding parameters for first bean if IsFirstBean is true
	--- and for second bean if IsFirstBean is false
	---


    Perform(me: in out);
    	---Purpose: 
    	--- Launches the algorithm
	--- 

    IsDone(me) returns Boolean from Standard;
    	---C++: inline
	---Purpose: 
    	--- Returns true if the computations was successfull
	--- otherwise returns false

    Result(me)
	returns SequenceOfRanges from XIntTools;
	---C++: return const &

    Result(me; theResults: out SequenceOfRanges from XIntTools);


    -- private

    ComputeRoughIntersection(me: in out)
    	is private;

    FastComputeIntersection(me: in out)
    	returns Boolean from Standard is private;
    
    ComputeUsingExtrema(me: in out; theRange2: Range from XIntTools)
    	is private;
    
    ComputeNearRangeBoundaries(me: in out; theRange2: Range from XIntTools)
    	is private;
    
    ComputeRangeFromStartPoint(me: in out; ToIncreaseParameter : Boolean from Standard;
    	    	   			   theParameter        : Real from Standard;
					   theIndex            : Integer from Standard;
					   theParameter2       : Real from Standard;
    	    	    	    	    	   theRange2           : Range from XIntTools)
    	is private;

    Distance(me: in out; theArg           : Real from Standard;
    	    	    	 theArgOnOtherBean: out Real from Standard)
    	returns Real from Standard
    	is private;

fields

    -- sources    
    myCurve1          : Curve   from BRepAdaptor;
    myCurve2          : Curve   from BRepAdaptor;
    myTrsfCurve1      : Curve from Geom;
    myTrsfCurve2      : Curve from Geom;

    myFirstParameter1 : Real from Standard;
    myLastParameter1  : Real from Standard;
    myFirstParameter2 : Real from Standard;
    myLastParameter2  : Real from Standard;

    myBeanTolerance1  : Real from Standard;
    myBeanTolerance2  : Real from Standard;
    
    myCurveResolution1: Real from Standard;
    myCriteria        : Real from Standard;

    -- tools
    myProjector      : ProjectPointOnCurve from GeomAPI;
    myRangeManager   : MarkedRangeSet from XIntTools;    
    myDeflection     : Real from Standard;

    -- results
    myResults        : SequenceOfRanges from XIntTools;

    myIsDone         : Boolean from Standard;

end BeanBeanIntersector from XIntTools;
