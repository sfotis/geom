-- Created on: 2001-12-13
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class PntOnFace from XIntTools 

	---Purpose: Contains a Face, a 3d point, corresponded UV parameters and a flag

uses
    Face from TopoDS, 
    Pnt  from  gp
--raises

is 
    Create 
    	returns PntOnFace from XIntTools;  
	---Purpose:
	--- Empty constructor
	---

    Init(me:out;  
    	 aF: Face from TopoDS; 
	 aP: Pnt  from  gp; 
	 U : Real from  Standard;     
	 V : Real from  Standard); 
	---Purpose:
	--- Initializes me by aFace, a 3d point
	--- and it's UV parameters on face
	---
	
    SetFace(me:out; 
    	    aF:Face from TopoDS); 
	---Purpose:
	--- Modifier
	---
	
    SetPnt (me:out; 
    	    aP:Pnt  from  gp);
    	---Purpose:
	--- Modifier
	---

    SetParameters (me:out; 
	    	   U : Real from  Standard;     
	    	   V : Real from  Standard);
    	---Purpose:
	--- Modifier
	---
	
    SetValid(me:out; 
	     bF : Boolean from Standard); 
    	---Purpose:
	--- Modifier
	---
	    	 
    Valid(me) 
	returns Boolean from Standard; 
	---Purpose:
	--- Selector
	---
	 
    Face(me) 
    	returns Face from TopoDS; 
    	---C++:  return const & 
	---Purpose:
	--- Selector
	---
     
    Pnt (me) 
    	returns Pnt  from gp; 
    	---C++:  return const & 
	---Purpose:
	--- Selector
	---

    Parameters (me; 
	    	U :out Real from Standard;     
	    	V :out Real from Standard); 
    	---Purpose:
	--- Selector
	---
	  
    IsValid(me) 
	returns Boolean from Standard; 
	---Purpose:
	--- Selector

fields  

    myIsValid : Boolean from Standard;    
    myPnt : Pnt  from  gp; 
    myU   : Real from  Standard;        
    myV   : Real from  Standard;        
    myFace: Face from TopoDS; 
end PntOnFace;
