-- Created on: 2002-02-04
-- Created by: Peter KURNEV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class WireShell from XBOP inherits WireShape from XBOP

	---Purpose: 
    	--  The class to perform a Boolean Operations (BO)       
	--  Common,Cut,Fuse  between arguments when one of them is  
    	--  a wire and other argument is a shell 
	--    	 
uses
    DSFiller  from XBOPTools, 
    PDSFiller from XBOPTools, 
    --modified by NIZHNY-MKK  Tue Sep  7 11:46:27 2004
    ShapeEnum from TopAbs,
    Operation from XBOP,
    ListOfShape from TopTools 
is
    Create   
    	returns  WireShell from XBOP; 
    	---Purpose:  
    	--- Empty constructor;
    	---
    Do  (me:out) 
    	is  redefined;  
    	---Purpose:  
    	--- See base classes, please 
    	---
    DoWithFiller      (me:out; 
    	     aDSF: DSFiller from XBOPTools) 
    	is  redefined; 
    	---Purpose:  
    	--- See base classes, please 
    	---
    Destroy (me: in out) 
    	is redefined; 
    	---C++: alias "Standard_EXPORT virtual ~XBOP_WireShell(){Destroy();}"  
    	---Purpose:  
    	--- Destructor 
    	---
    BuildResult (me:out) 
	is  redefined;	 
    	---Purpose:  
    	--- See base classes, please 
    	---
    --modified by NIZHNY-MKK  Tue Sep  7 11:46:00 2004
    CheckArgTypes(myclass; theType1, theType2: ShapeEnum from TopAbs;
    	    	    	   theOperation: Operation from XBOP) 
	 returns Boolean from Standard;  
    	---Purpose: 
    	--- Check the types of arguments.      
    	--- Returns  FALSE if types of arguments     
    	--- are non-valid to be  treated by the         
    	--- agorithm
    
    CheckArgTypes(me) 
	returns Boolean from Standard 
    	is  private;  
    	---Purpose:  
    	--- Internal  usage
    	---
    
--fields

end WireShell;
