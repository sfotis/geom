-- Created on: 2000-05-22
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Root from XIntTools 

	---Purpose: The class is to describe the root of  
        --          function of one variable  for  Edge/Edge 
	--          and  Edge/Surface  algorithms. 
	
uses 
    State  from  TopAbs

---raises
is 
    Create  
    	returns Root from XIntTools ; 
    	---Purpose: 
    	--- Empty constructor
	---
     
    Create(aRoot:  Real    from Standard; 
    	   aType:  Integer from Standard) 
    	returns Root from XIntTools ;  
    	---Purpose: 
	--- Initializes my by range of parameters
	--- and type of root
	---
	    		  
    SetRoot  (me:out;  aRoot:  Real from Standard); 
    	---Purpose: 
    	--- Sets the Root's value
	---
   
    SetType  (me:out;  aType:  Integer from Standard); 
    	---Purpose: 
    	--- Sets the Root's Type
	---
    
    SetStateBefore  (me:out;  aState: State  from  TopAbs); 
    	---Purpose: 
    	--- Set  the  value of the state before the root   
    	--- (at  t=Root-dt)
	---

    SetStateAfter   (me:out;  aState: State  from  TopAbs); 
    	---Purpose: 
    	--- Set  the  value of the state after the root   
    	--- (at  t=Root-dt)
	---

    SetLayerHeight  (me:out;  aHeight:Real from Standard); 
    	---Purpose: 
    	--- Not  used  in  Edge/Edge  algorithm 
	---

    SetInterval     (me:out;  t1, t2, f1, f2:Real from Standard); 
    	---Purpose: 
    	--- Sets the  interval  from which the Root was 
    	--- found [t1,t2] and the  corresponding  values   
    	--- of  the  function  on  the  bounds f(t1), f(t2).
	---
     
    Root  (me)   
    	returns Real from Standard; 
    	---Purpose: 
    	--- Returns the Root  value 
	---
     
    Type  (me)       
      	returns Integer from Standard;  
    	---Purpose: 
    	--- Returns the  type  of  the  root 
    	--- =0  -  Simple (was  found  by  bisection  method); 
    	--- =2  -  Smart when f1=0, f2!=0 or  vice  versa 
    	---        (was  found  by  Fibbonacci method); 
    	--- =1  -  Pure   (pure  zero  for all t [t1,t2] ); 
    
    StateBefore(me) 
    	returns State  from  TopAbs;
    	---Purpose: 
    	--- Returns the state before the root
	---

    StateAfter(me) 
    	returns State  from  TopAbs;  
    	---Purpose: 
    	--- Returns the state after the root
	---

    LayerHeight (me) 
	returns Real from Standard;  
    	---Purpose: 
    	--- Not  used  in  Edge/Edge  algorithm
	---

    IsValid   (me) 
    	returns  Boolean  from Standard; 
    	---Purpose: 
    	--- Returns the validity flag for the root, 
    	--- True if   
    	--- myStateBefore==TopAbs_OUT && myStateAfter==TopAbs_IN or	     
    	--- myStateBefore==TopAbs_OUT && myStateAfter==TopAbs_ON or	     
    	--- myStateBefore==TopAbs_ON  && myStateAfter==TopAbs_OUT or 
    	--- myStateBefore==TopAbs_IN  && myStateAfter==TopAbs_OUT  . 
    	--- For  other  cases it  returns  False. 
	---
     
    Interval  (me;  t1:out Real from Standard;  
    	    	    t2:out Real from Standard;  
    	    	    f1:out Real from Standard;  
    	    	    f2:out Real from Standard); 
    	---Purpose: 
    	--- Returns the values of interval  from which the Root was 
    	--- found [t1,t2] and the  corresponding  values   
    	--- of  the  function  on  the  bounds f(t1), f(t2).
	---

fields 
    myRoot:  Real from Standard;
    
    myType:  Integer from Standard; 
     
    myLayerHeight:  Real from Standard;
    myStateBefore:  State  from  TopAbs; 
    myStateAfter :  State  from  TopAbs; 

    myt1:  Real from Standard;
    myt2:  Real from Standard;
    myf1:  Real from Standard;
    myf2:  Real from Standard;
end Root;
