-- Created on: 1996-01-05
-- Created by: Jean Yves LEBEY
-- Copyright (c) 1996-1999 Matra Datavision
-- Copyright (c) 1999-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


deferred class CompositeClassifier from XBOP inherits LoopClassifier from XBOP

    ---Purpose:  
    --  The Root class for algorithms  
    --  to   classify composite Loops, i.e, Loops that  
    --  can be either a Shape, or a block of Elements.
    --   
    
uses
    
    ShapeEnum from TopAbs,
    Shape     from TopoDS,
    State     from TopAbs,
     
    Loop         from XBOP,
    BlockBuilder from XBOP
    
is

    Initialize(BB : BlockBuilder from XBOP);
    	---Purpose:  
    	--- Initializing the object with BlockBuilder;   
    	---
    Compare(me :out;  
    	L1 : Loop from XBOP;  
    	L2 : Loop from XBOP)  
    	returns State from TopAbs
    	is redefined;
    	---Purpose:  
    	--- Classify loop <L1> with  <L2>  
    	---
    CompareShapes(me :out;  
    	B1 : Shape from TopoDS;
    	B2 : Shape from TopoDS)
    	---Purpose:  
    	--- Classify shape <B1> with shape <B2>
    	---
	returns State from TopAbs  
    	is deferred;
    
    CompareElementToShape(me :out;  
    	E : Shape from TopoDS;
    	B : Shape from TopoDS) 
    	returns State from TopAbs  
    	is deferred;
    	---Purpose:  
    	--- Classify element <E> with shape <B>
    	---
    ResetShape(me :out;  
    	B : Shape from TopoDS)  
    	is deferred;
    	---Purpose:  
    	--- Prepare classification involving shape <B>
    	--- Calls ResetElement on first element of <B>
	---
    
    ResetElement(me :out;  
    	E : Shape from TopoDS)  
    	is deferred;
    	---Purpose:  
    	--- Prepare classification involving element <E>.
    	---
    CompareElement(me :out;  
    	E : Shape from TopoDS)  
    	is deferred;
    	---Purpose:  
    	--- Add element <E> in the set of elements used in classification.
    	---
    State(me :out)  
    	returns State from TopAbs  
    	is deferred;
    	---Purpose:  
    	--- Returns state of classification of 2D point, defined by 
    	--- ResetElement, with the current set of elements,  
    	--- defined by Compare.
    	---
fields

    myBlockBuilder : Address  
    	is protected; 

end CompositeClassifier;
