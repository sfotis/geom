-- Created on: 2001-05-18
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Section from XBOP inherits Builder from XBOP

	----Purpose: Performs the Boolean Operation (BO) Section 
    	---          for the shapes   
	

uses
    DSFiller from XBOPTools,
    HistoryCollector from XBOP

is
    Create 
    	returns Section from XBOP; 
    	---Purpose:  
    	--- Empty constructor;  
    	---
    Do  (me:out) 
    	is  redefined;
    	---Purpose: 
    	--- Does the BO from the beggining to the end, 
    	--- i.e.  create new DataStructure, DSFiller,         
    	--- compute all  interferences, compute states, 
    	--- build result etc 
    	---
    Do  (me:out;toApprox         : Boolean from Standard;
    	    	toComputePCurve1 : Boolean from Standard;
    	    	toComputePCurve2 : Boolean from Standard);
    	---Purpose: 
    	--- Does the BO from the beggining to the end, 
    	--- i.e.  create new DataStructure, DSFiller,         
    	--- compute all  interferences, compute states, 
    	--- build result etc 
    	---

    DoWithFiller (me:out; 
    	    	  aDSF: DSFiller from XBOPTools) 
    	is  redefined; 
    	---Purpose:   
    	--- Does the BO using existing Filler to the end        
    	---
      
    Destroy (me: in out) 
    	is redefined; 
    	---C++: alias "Standard_EXPORT virtual ~XBOP_Section(){Destroy();}"   	 
    	---Purpose:    
    	--- Destructor 
    	---

    SetHistoryCollector(me: in out; theHistory: HistoryCollector from XBOP)
    	is redefined virtual;

--fields 

end Section;
