-- Created on: 2001-04-09
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class ShellSplitter from XBOP 

	---Purpose:  
    	---  the algorithm to split (multiconnexed)   
    	---  shells on a solid onto biconnexed shells 
	---  when each edge is shared by only two or one  
    	--   faces       

uses 

    Shell  from TopoDS,
    ListOfShape from  TopTools, 
    
    ListOfListOfShape from XBOPTColStd, 
    
    EdgeInfo                         from XBOP,
    IndexedDataMapOfEdgeListFaceInfo from XBOP

 --raises

is 
    Create   
    	returns ShellSplitter from XBOP; 
    	---Purpose:  
    	--- Empty constructor; 
    	---
    DoWithListOfEdges(me:out; 
    	    	aLE:ListOfShape from  TopTools); 
    	---Purpose:  
    	--- Perform the algorithm using the  list of shapes <aLE> as data  
    	---
    SetShell    (me:out; 
		aShell:Shell from TopoDS);    	     
    	---Purpose:  
    	--- Modifier
    	---
    Shell    (me) 
	returns Shell from TopoDS; 
    	---C++:  return const &	 
    	---Purpose:  
    	--- Selector
    	---
    DoWithShell (me:out); 
    	---Purpose:  
    	--- Perform the algorithm using the shell as data  
    	---
    Do          (me:out) 
    	is private;  
    	---Purpose:  
    	--- Perform the algorithm 
    	---
    IsNothingToDo (me) 
    	returns  Boolean from Standard;
    	---Purpose: 
    	--- Returns TRUE if the source shell is valid and      
    	--- there  is  nothing to correct 
    	---
    IsDone (me) 
    	returns  Boolean from Standard; 
    	---Purpose:  
    	--- Returns TRUE if the algorithm was performed  
    	--- successfuly 
	---
    Shapes (me) 
    	returns  ListOfListOfShape from XBOPTColStd;
    	---C++:  return const &	    		 
    	---Purpose:  
    	--- Selector
    	---
    
	
fields  
    myShell      :  Shell from TopoDS;
    myIsDone     :  Boolean from Standard;
    myNothingToDo:  Boolean from Standard;
    myShapes     :  ListOfListOfShape from XBOPTColStd; 
    mySmartMap   :  IndexedDataMapOfEdgeListFaceInfo from XBOP;  
    myFaces      :  ListOfShape from  TopTools; 
    
end ShellSplitter;










