-- Created on: 2001-02-08
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class Pave from XBOPTools 

	---Purpose:  
    	--  Class for storing info about a vertex on an edge 

uses 
    KindOfInterference from XBooleanOperations 
    
is 
    Create 
    	returns Pave from XBOPTools; 
    	---Purpose:  
    	--- Empty constructor 
    	---
    Create (Index: Integer from Standard; 
            aParam:Real from Standard;  
    	    aType:  KindOfInterference from XBooleanOperations   
    	    	    =XBooleanOperations_UnknownInterference)   
    	returns Pave from XBOPTools;  
    	---Purpose:  
    	--- Constructor 
    	--- Index  - DS-index of the vertex    	 
    	--- aParam - value of the parameter of the vertex on an edge              
    	--- aType  - the type of interference from which the pave comes from        
    	---
    SetParam  (me:out; aParam:Real from Standard);  
    	---Purpose:  
    	--- Modifier  
    	---
    SetIndex  (me:out; Index: Integer from Standard); 
    	---Purpose:  
    	--- Modifier  
    	---
    SetType   (me:out;  aType:KindOfInterference from XBooleanOperations); 
    	---Purpose:  
    	--- Modifier  
    	---
    SetInterference (me:out; Index: Integer from Standard); 
    	---Purpose:  
    	--- Modifier  
    	--- Sets the index of the interference in corresponding table 
    	---
    Param     (me) 
    	returns Real from Standard;	    		  
    	---Purpose:  
    	--- Selector  
    	---
    Index     (me) 
	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector  
    	---
    Type   (me) 
    	returns KindOfInterference from XBooleanOperations; 
    	---Purpose:  
    	--- Selector  
    	---
    Interference(me) 
	returns Integer from Standard; 
    	---Purpose:  
    	--- Selector  
    	---
    IsEqual(me;  Other:Pave from XBOPTools) 
    	returns Boolean from Standard; 
    	---Purpose:  
    	--- Returns TRUE if  <Other>==me 
    	---
fields 
    myParam:  Real from Standard; 
    myIndex:  Integer from Standard; 
    myType :  KindOfInterference from XBooleanOperations; 
    myInterf: Integer from Standard; 
end Pave;


