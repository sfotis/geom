-- Created on: 2001-04-09
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class WireSplitter from XBOP 

    	---Purpose: 
    	---  the algorithm to split multiconnexed   
    	---  wires on a face onto biconnexed ones 
	---  .
uses
    Face   from TopoDS,  
    Vertex from TopoDS, 
    Edge   from TopoDS, 
    
    SequenceOfPnt2d  from TColgp, 
    SequenceOfShape  from TopTools,   
    ListOfShape      from TopTools, 
    
    ListOfListOfShape from XBOPTColStd, 
    
    EdgeInfo                           from XBOP,
    IndexedDataMapOfVertexListEdgeInfo from XBOP

--raises

is 
    Create   
    	returns WireSplitter from XBOP; 
    	---C++: inline
    	---Purpose:  
    	--- Empty constructor; 
    	---
    SetFace  (me:out; 
    	    	aF: Face from TopoDS); 
    	---C++: inline
    	---Purpose:  
    	--- Modifier
    	---
    DoWithListOfEdges(me:out; 
    	    	    	aLE:ListOfShape from  TopTools); 
    	---Purpose:  
    	--- Perform the algorithm using the  list of shapes <aLE> as data  
    	---
    DoWithFace  (me:out); 
    	---Purpose:  
    	--- Perform the algorithm using the face as data  
    	---
    Do          (me:out) 
    	is private;  
    	---Purpose:  
    	--- Perform the algorithm 
    	---
    IsNothingToDo (me) 
    	returns  Boolean from Standard;
    	---C++: inline
    	---Purpose:  
    	--- Returns TRUE if the source wire is biconnexed and      
    	--- there is nothing to correct 
    	---
    IsDone (me) 
    	returns  Boolean from Standard; 
    	---C++: inline
    	---Purpose:  
    	--- Returns TRUE if the algorithm was performed  
    	--- successfuly
	---
    Face   (me) 
    	returns Face from TopoDS; 
    	---C++:  return const &	    	 
    	---C++: inline
    	---Purpose:  
    	--- Selector
    	---
    Shapes (me) 
    	returns  ListOfListOfShape from XBOPTColStd; 
    	---C++:  return const &	    		 
    	---C++: inline
    	---Purpose:  
    	--- Selector
    	---
    
	
fields  

    myFace       :  Face from TopoDS; 
    myIsDone     :  Boolean from Standard;
    myNothingToDo:  Boolean from Standard;
    myShapes     :  ListOfListOfShape from XBOPTColStd; 
    mySmartMap   :  IndexedDataMapOfVertexListEdgeInfo from XBOP;  
    myEdges      :  ListOfShape from  TopTools; 
    
end WireSplitter;
