-- Created on: 2002-02-01
-- Created by: Peter KURNEV
-- Copyright (c) 2002-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class WireWire from XBOP inherits WireShape from XBOP

	---Purpose: 
    	---        
    	---        Performs Boolean Operations  (BO)  
    	---        Common,Cut,Fuse for wires as      
	---        arguments 
uses
    DSFiller  from XBOPTools, 
    PDSFiller from XBOPTools, 
    ListOfShape from TopTools 
    
--raises

is 
    Create   
    	returns  WireWire from XBOP; 
    	---Purpose:  
    	--- Empty constructor;
    	---
    Do  (me:out) 
    	is  redefined; 	 
    	---Purpose:  
    	--- (See base classes, please)
    	---
    DoWithFiller      (me:out; 
    	     aDSF: DSFiller from XBOPTools) 
    	is  redefined; 
    	---Purpose:  
    	--- (See base classes, please)
    	---
    Destroy (me: in out) 
    	is redefined; 
    	---C++: alias "Standard_EXPORT virtual ~XBOP_WireWire(){Destroy();}"  
    	---Purpose:   
    	--- Destructor 
    	---
    BuildResult (me:out) 
	is  redefined;	 
    	---Purpose:  
    	--- See base classes, please 
    	---
    
--fields
  
end WireWire;
