-- Created on: 2001-06-25
-- Created by: Michael KLOKOV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.


class ShellFaceClassifier from XBOP inherits CompositeClassifier from XBOP


    	---Purpose:  
	
    	--- The  algorithm is to classify loops that  
    	--  consist of faces and shells
	--- 
    
uses
    
    Shape               from TopoDS,
    Shell               from TopoDS,
    State               from TopAbs,
    Pnt                 from gp,
    Builder             from BRep, 
    BlockBuilder        from XBOP,
    SolidClassifier     from XBOP,
    DataMapOfShapeShape from TopTools

is
    Create(theBlockBuilder: BlockBuilder from XBOP)
    	returns ShellFaceClassifier from XBOP;
    	---Purpose: 
    	--- Creates a classifier in 3D space, to compare
    	--- a face with a set of faces,
    	--- a shell with a set of faces,
    	--- a shell with a shell
    	---
    Clear(me: in out);
    	---Purpose:  
    	--- Clears  contents of internal state of the object     
    	---
    CompareShapes(me : in out;  
    	    	  B1 : Shape from TopoDS;  
    	    	  B2 : Shape from TopoDS)
    	returns State from TopAbs
    	is redefined;
    	---Purpose:  
    	--- Classify shape <B1> with shape <B2> 
    	---
    CompareElementToShape(me : in out;  
    	    	  E : Shape from TopoDS;  
    	    	  B : Shape from TopoDS)
    
    	returns State from TopAbs
	is redefined;
    	---Purpose:  
    	--- Classify element <E> with shape <B> 
    	---
    ResetShape(me : in out;  
    	          B : Shape from TopoDS)
    	is redefined;
    	---Purpose:  
    	--- Prepare classification involving shape <B>
    	--- Calls ResetElement on first element of <B> 
    	---
    ResetElement(me : in out;  
    	          E : Shape from TopoDS)
	is redefined;
    	---Purpose:  
    	--- Prepare classification involving element <E>. 
    	---
    CompareElement(me : in out;  
    	    	  E : Shape from TopoDS);
    	---Purpose:  
    	--- Add element <E> in the set of elements used in classification.
    	---
    State(me : in out)  
    	returns State from TopAbs
	is redefined;
    	---Purpose:  
    	--- Returns state of classification of 2D point, defined by 
    	--- ResetElement, with the current set of elements,  
    	--- defined by Compare. 
    	---
    
fields

    myFirstCompare:    Boolean from Standard;
    myPoint:           Pnt from gp;
    myShell:           Shell from TopoDS;
    myBuilder:         Builder from BRep;
    mySolidClassifier: SolidClassifier from XBOP; 
    myFaceShellMap :   DataMapOfShapeShape from TopTools;

end ShellFaceClassifier from XBOP;
