-- Created on: 2000-11-21
-- Created by: Peter KURNEV
-- Copyright (c) 2000-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SSInterference from XBOPTools  
    inherits ShapeShapeInterference from XBOPTools 

	---Purpose: class for storing a Face/Face interference     
	---         Each  F/F interference  contains  information  about 
	---         1.  myPBs   - PaveBlocks (made from edges from the faces  
    	---             that are IN-2D or ON-2D;    
	---         2.  myCurves- Sequence of curves of intersection;      
	---         3.  myTangentFacesFlag  - The BOOL flag indicates that  
	---             the  faces are SD in terms of the F/F Intersector.     
	---         4.  mySenseFlag  - value that is equal +1 or -1 depending 
	---             on scalar product between normals to each face.  This      
	---             valie is valid for the SDF only.        
	---         5.  myAlonePnts  - contains 3D-points that are place 
	---             of  intersection between the two faces    
        ---         6.  myAloneVertices   - contains indices of vertices  
	---             that correspond to the points  myAlonePnts; 
	---

uses   

    PaveBlock        from XBOPTools, 
    PaveSet          from XBOPTools,
    ListOfPaveBlock  from XBOPTools, 
    SequenceOfCurves from XBOPTools, 
    IndexedDataMapOfIntegerState from XBOPTools, 

    SequenceOfCurves      from XIntTools,  
    SequenceOfPntOn2Faces from XIntTools, 

    ListOfInteger from  TColStd    
    --
is 
    Create  
    	returns  SSInterference from XBOPTools; 
    	---Purpose:  
    	--- Empty constructor  
    	---
    Create  (anIndex1: Integer  from Standard;
    	     anIndex2: Integer  from Standard; 
    	     aTolR3D : Real from Standard; 
    	     aTolR2D : Real from Standard; 
    	     aCurves : SequenceOfCurves from XIntTools; 
    	     aPnts   : SequenceOfPntOn2Faces from XIntTools) 	
    	returns SSInterference from XBOPTools;  
    	---Purpose:   
    	--- Constructor 
    	--- anIndex1,  
    	--- anIndex2 see XBOPTools_ShapeShapeInterference for details     
    	--- aTolR3D  - value of tolerance to reach in 3D-space      
    	--- aTolR2D  - value of tolerance to reach in 2D-space      
    	--- aCurves  see  XIntTools_Curve  for details,  please 
    	---
    AppendBlock(me:out;   
    	    	aPB:PaveBlock from XBOPTools);      
    	---Purpose:  
    	--- Modifier 
    	---
    PaveBlocks(me) 
    	returns ListOfPaveBlock from XBOPTools; 
    	---C++:  return const & 
    	---Purpose:  
    	--- Selector  
    	---
    NewPaveSet(me:out) 
    	returns PaveSet from XBOPTools; 
    	---C++:  return &	 
    	---Purpose:  
    	--- Selector  
    	---
    TolR3D  (me) 
    	returns Real from Standard;            
    	---Purpose:  
    	--- Selector  
    	---
    TolR2D  (me) 
    	returns Real from Standard;
    	---Purpose:  
    	--- Selector  
    	---
    Curves(me:out) 
    	returns SequenceOfCurves from XBOPTools; 
    	---C++:  return &   
    	---Purpose:  
    	--- Selector  
    	---
    SetTangentFacesFlag(me:out; 
    	    aFlag:Boolean from Standard); 
    	---Purpose:  
    	--- Modifier  
    	---
    IsTangentFaces(me) 
    	returns Boolean from Standard; 
    	---Purpose:  
    	--- Selector  
    	---
    SetSenseFlag (me:out;  
    	aFlag:Integer from Standard);      
    	---Purpose:  
    	--- Modifier  
    	---
    SenseFlag (me)  
    	returns Integer from Standard; 	 
    	---Purpose:  
    	--- Selector  
    	---
    SetStatesMap(me:out; 
    	aStatesMap:  IndexedDataMapOfIntegerState from XBOPTools); 
    	---Purpose: 
    	--- Modifier  
    	---
    StatesMap(me)  
    	returns  IndexedDataMapOfIntegerState from XBOPTools;  
    	---C++:  return const &  	
    	---Purpose: 
    	--- Selector  
    	---
    SetAlonePnts(me:out;  
    	aPnts:SequenceOfPntOn2Faces from XIntTools); 
    	---Purpose:  
    	--- Modifier  
    	---
    AlonePnts(me) 
    	returns SequenceOfPntOn2Faces from XIntTools; 
    	---C++:  return const &  	 
    	---Purpose:  
    	--- Selector
    	---
    AloneVertices(me:out) 
    	returns ListOfInteger from  TColStd; 
    	---C++:  return &  
    	---Purpose:  
    	--- Selector 
    	---  
    --modified by NIZNHY-PKV Fri Jun 30 10:05:36 2006f	
    SetSharedEdges(me:out;  	 
	    aLS:ListOfInteger from TColStd); 
        ---Purpose:  
    	--- Modifier  
    	---    
    SharedEdges(me)  	 
	returns ListOfInteger from TColStd;  
    	---C++:  return const &  
    	---Purpose:  
    	--- Selector 
    	---      
    --modified by NIZNHY-PKV Fri Jun 30 10:05:41 2006t 
     
fields
    
    myPBs         : ListOfPaveBlock from XBOPTools is protected;  
    myNewPaveSet  : PaveSet from XBOPTools is protected;
    myTolR3D      : Real from Standard is protected; 
    myTolR2D      : Real from Standard is protected; 
     
    myCurves           : SequenceOfCurves from XBOPTools is protected;  
    myAlonePnts        : SequenceOfPntOn2Faces from XIntTools is protected; 
    myAloneVertices    : ListOfInteger from  TColStd is protected; 

    myTangentFacesFlag : Boolean from Standard is protected; 
    mySenseFlag        : Integer from Standard is protected;  	     
    myStatesMap        : IndexedDataMapOfIntegerState from XBOPTools is protected;
--modified by NIZNHY-PKV Fri Jun 30 10:02:27 2006f   
    mySharedEdges      : ListOfInteger from TColStd is protected;   
--modified by NIZNHY-PKV Fri Jun 30 10:02:34 2006     
end SSInterference;
