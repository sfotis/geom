-- Created on: 2001-06-06
-- Created by: Peter KURNEV
-- Copyright (c) 2001-2012 OPEN CASCADE SAS
--
-- The content of this file is subject to the Open CASCADE Technology Public
-- License Version 6.5 (the "License"). You may not use the content of this file
-- except in compliance with the License. Please obtain a copy of the License
-- at http://www.opencascade.org and read it completely before using this file.
--
-- The Initial Developer of the Original Code is Open CASCADE S.A.S., having its
-- main offices at: 1, place des Freres Montgolfier, 78280 Guyancourt, France.
--
-- The Original Code and all software distributed under the License is
-- distributed on an "AS IS" basis, without warranty of any kind, and the
-- Initial Developer hereby disclaims all such warranties, including without
-- limitation, any warranties of merchantability, fitness for a particular
-- purpose or non-infringement. Please see the License for the specific terms
-- and conditions governing the rights and limitations under the License.



class SDFWESFiller from XBOP 

	---Purpose:  
    	--  The  algorithm that fills a wire edges set (WES) 
    	--  for a couple of faces that are same domain 
    	--- 
	
uses 
    Face from TopoDS, 
    ListOfShape from TopTools,
    DSFiller  from XBOPTools, 
    PDSFiller from XBOPTools, 
    IndexedDataMapOfIntegerState from XBOPTools,  
    
    Operation    from XBOP,  
    WireEdgeSet  from XBOP,
    PWireEdgeSet from XBOP 
    
    
--raises

is 
    Create   
    	returns SDFWESFiller from XBOP; 
    	---Purpose:  
    	--- Empty constructor
    	---
    Create  (nF1: Integer from Standard; 
    	     nF2: Integer from Standard; 
    	     aDSF: DSFiller from XBOPTools);
    	---Purpose:  
    	--- Constructor
    	--- nF1, nF2 - indices of faces in the DataStructue (DS)    
    	---
    SetStatesMap(me:out; 
    	aStatesMap:  IndexedDataMapOfIntegerState from XBOPTools); 
    	---Purpose: 
    	--- Modifier  
    	---
    SetFaces(me:out; 
    	nF1: Integer from Standard;  
    	nF2: Integer from Standard);  
    	---Purpose: 
    	--- Modifier  
    	---
    SetDSFiller(me:out; 
    	aDSF: DSFiller from XBOPTools); 
    	---Purpose: 
    	--- Modifier  
    	---
    SetOperation (me:out; 
    	    	  anOp:Operation from XBOP);   
    	---Purpose: 
    	--- Modifier  
    	---
    SetSenseFlag (me:out;  
    	aFlag:Integer from Standard); 
    	---Purpose: 
    	--- Modifier 
    	--- Assigns sensitivity flag for the faces in accordance 
    	--- with scalar product between theirs normalls 
    	--- 1  for same sense;  -1 for different sense      
    	---

    Prepare(me:out); 
    	---Purpose: 
    	--- Prepares data for the algorithm 
    	---
    Do  (me:out; 
    	 aWES:WireEdgeSet from XBOP); 
    	---Purpose:  
    	--- Performs the algorithm 
    	---
    DSFiller(me) 
    	returns DSFiller from XBOPTools; 
    	---C++:  return const & 
    	---Purpose: 
    	--- Selector  
    	---
    StatesMap(me)  
    	returns  IndexedDataMapOfIntegerState from XBOPTools;  
    	---C++:  return const &  	
    	---Purpose: 
    	--- Selector  
    	---
    Faces(me; 
    	nF1:out Integer from Standard;  
    	nF2:out Integer from Standard); 
    	---Purpose: 
    	--- Selector  
    	---
    SenseFlag (me)  
    	returns Integer from Standard; 	     
    	---Purpose: 
    	--- Selector  
    	---
    Operation  (me) 
    	returns Operation from XBOP; 
    	---Purpose: 
    	--- Selector  
    	---
    AssignStates (me:out;      
    	    	    nF1: Integer from Standard;  
    	    	    nF2: Integer from Standard) 
    	is  private;  
    	---Purpose: 
    	--- Assigns the 2D-State for split parts of  
    	--- the edges having 3D-Curves of given faces       	     
    	--- Internal  Purpose
    	---
    PrepareOnParts(me:out) 
    	is  private;  
    	---Purpose: 
    	--- Prepares ON 2D parts to filled the WES  
    	--- Internal Purpose 
    	---
    PrepareWESForZone(me:out;      
    	    	    nF1: Integer from Standard;  
    	    	    nF2: Integer from Standard) 
    	is  private;
    	---Purpose: 
    	--- Fills the WES by split parts of the edges for         
    	--- the Common Zone  
    	--- Internal Purpose 
    	---
    PrepareWESForCut(me:out;      
    	    	    nF1: Integer from Standard;  
    	    	    nF2: Integer from Standard) 
    	is  private;
    	---Purpose: 
    	--- Fills the WES by split parts of the edges for         
    	--- the Cut operation 
    	--- Internal Purpose 
    	--- 
    PrepareOnParts(me:out; 
    	    	    nF1: Integer from Standard;  
    		    nF2: Integer from Standard; 
    	    	    Op : Operation from XBOP) 
    	is  private; 
    	---Purpose: 
    	--- Fills the WES by split parts (ON 2D) of the edges 
    	--- Internal Purpose  
    	---
    PrepareFaces(me; 
		   nF1: Integer from Standard;  
    		   nF2: Integer from Standard;  
		   aF1:out Face from TopoDS;
		   aF2:out Face from TopoDS) 
    	is  private;
    	---Purpose: 
    	--- Make orientation of the faces consistent  
    	--- Internal Purpose 
    	---
    AssignDEStates (me:out; 
    	    	    nF1: Integer from Standard;  
    		    nF2: Integer from Standard) 
    	is  private; 
    	---Purpose:  
    	--- Assigns the 2D-State for split parts of  
    	--- the edges that do not have 3D-Curves of given faces   
    	--- Internal Purpose 
    	---
    AssignDEStates (me:out; 
    	    	    nF1: Integer from Standard;  
    		    nE1: Integer from Standard; 
    		    nF2: Integer from Standard) 
    	is  private; 
    	---Purpose: 
    	--- Assigns the 2D-State for split parts of  
    	--- the edge  nE1 that do not have 3D-Curves from face nF1 
    	---
    	--- Internal Purpose 
    	---
    UpdateDEStates3D  (me:out); 
    	---Purpose:	 
    	--- Update 3D-State for edges    
    	---
    RejectedOnParts(me) 
    	returns ListOfShape from TopTools; 
    ---C++: return const &   
    ---Purpose:   
    --  Returns all split edges of nF1 that are CB with 
    --  splis of nF1 but not included in myWES,     
    
fields
 
    myDSFiller  : PDSFiller from XBOPTools; 
    myOperation : Operation from XBOP;
    myNF1       : Integer from Standard; 
    myNF2       : Integer from Standard; 
      
    myWES       : PWireEdgeSet from XBOP; 
    myStatesMap:  IndexedDataMapOfIntegerState from XBOPTools;
    mySenseFlag:  Integer from Standard;   
    myRejectedOnParts: ListOfShape  from TopTools;  
     
end SDFWESFiller;

